module Menu_Pixel_Gen ();
    
endmodule