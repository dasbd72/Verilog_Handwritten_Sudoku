/*
    clk : posedge clock signal
    rst : posedge reset signal
    start : req 1 cycle signal
    layer_input : req 784 cycle
    layer_0 : last until next start signal
    finish : last 1 cycle
 */
module Dense_0(
    input  wire clk, 
    input  wire rst,
    input  wire start,
    input  wire [28*28 - 1:0] layer_input,
    output reg  [16*64 - 1:0] layer_0,
    output reg  finish
    );
    localparam HEIGHT = 784;
    localparam WIDTH = 64;
    localparam [802815:0] kernel_0 = {16'h001a,16'h002a,-16'h0017,-16'h004e,16'h0013,16'h0000,-16'h001e,16'h0037,16'h0059,-16'h0021,-16'h000c,16'h0021,16'h0013,16'h005b,-16'h0016,-16'h005e,-16'h002c,16'h003f,-16'h000c,16'h001c,-16'h002d,16'h0063,-16'h0004,16'h000a,-16'h0004,16'h0003,-16'h002a,-16'h0005,-16'h000d,-16'h0001,-16'h0043,-16'h0026,-16'h0012,-16'h004f,-16'h003e,-16'h002f,-16'h0049,-16'h002b,16'h0070,-16'h003c,-16'h0023,16'h0054,-16'h0001,16'h0081,16'h0024,16'h002f,-16'h0037,-16'h002a,16'h007f,16'h0010,16'h003a,-16'h0027,-16'h001b,-16'h0015,-16'h005e,16'h0018,16'h005a,-16'h0079,16'h0025,16'h0019,16'h0066,16'h000e,-16'h001a,-16'h004a,-16'h0016,16'h0011,-16'h001c,-16'h0037,16'h0044,16'h0014,16'h0010,16'h001a,16'h000b,-16'h005f,-16'h0002,-16'h0004,16'h0005,16'h0064,-16'h0011,-16'h007e,-16'h000f,16'h002c,-16'h002d,16'h000b,-16'h0009,16'h002f,16'h001d,-16'h0011,16'h0028,16'h0023,-16'h004b,16'h000a,16'h0016,16'h001b,-16'h002e,-16'h000a,-16'h0009,-16'h001e,-16'h0032,-16'h0021,-16'h0038,-16'h0009,16'h0092,16'h000c,-16'h0043,16'h0055,-16'h000d,16'h0059,16'h000b,16'h0039,-16'h0034,-16'h0022,16'h0086,16'h000c,16'h0029,-16'h0023,-16'h0029,-16'h0006,-16'h0019,16'h002f,16'h0047,-16'h0086,16'h0024,16'h000c,16'h0043,-16'h0002,-16'h0035,-16'h0041,-16'h0033,16'h000b,-16'h0048,-16'h0030,16'h002e,16'h0039,16'h0002,-16'h000a,16'h0014,-16'h007f,16'h0016,16'h0013,-16'h000e,16'h006b,-16'h0002,-16'h007e,-16'h0004,16'h0048,-16'h0047,16'h0022,-16'h0021,16'h0019,-16'h0011,-16'h0015,16'h003e,16'h0002,-16'h0053,16'h000b,16'h0014,16'h0003,-16'h0014,-16'h0013,16'h0010,-16'h0030,-16'h0013,-16'h0012,-16'h0056,16'h0016,16'h00a5,16'h0026,-16'h0044,16'h0048,-16'h001e,16'h0070,16'h002e,16'h003b,-16'h001b,-16'h000e,16'h0069,16'h000b,16'h0047,-16'h002b,-16'h002e,-16'h000b,-16'h0022,16'h0009,16'h0060,-16'h0050,16'h002e,16'h0013,16'h0015,16'h0010,-16'h005c,-16'h0059,-16'h002f,16'h0019,-16'h0072,-16'h001d,16'h002d,16'h004c,16'h0000,16'h0004,16'h0003,-16'h006d,16'h0017,-16'h000a,-16'h0025,16'h0073,16'h000c,-16'h0051,16'h0015,16'h0046,-16'h0060,16'h0011,16'h0000,16'h004c,16'h0012,-16'h0041,16'h0048,16'h0027,-16'h003f,16'h000c,16'h000d,16'h0010,-16'h0010,-16'h000c,16'h003d,-16'h001d,-16'h000c,16'h0001,-16'h007a,16'h0000,16'h00d8,16'h0015,-16'h0069,16'h0041,16'h0001,16'h0078,16'h003d,16'h006a,-16'h003c,-16'h0008,16'h006b,-16'h0019,16'h0046,-16'h003e,-16'h0068,-16'h000e,-16'h0034,-16'h0001,16'h003f,-16'h000a,16'h0021,16'h000b,-16'h001e,16'h0014,-16'h003e,-16'h0075,-16'h0051,16'h0033,-16'h007c,16'h0000,16'h006d,16'h0020,16'h0005,-16'h0011,-16'h0016,-16'h0050,16'h0004,-16'h002c,-16'h005a,16'h0055,-16'h0008,16'h0000,16'h0030,16'h0009,-16'h006d,16'h0002,16'h0000,16'h0044,16'h0012,-16'h006d,16'h003b,16'h002b,-16'h0028,16'h001e,16'h0020,16'h0005,-16'h001c,16'h000c,16'h002a,-16'h0013,-16'h0029,16'h0028,-16'h008d,16'h001a,16'h00d7,16'h000b,-16'h0061,16'h0050,16'h0007,16'h0060,16'h0014,16'h007f,-16'h0041,16'h0016,16'h006c,-16'h001d,16'h0035,-16'h005e,-16'h007e,-16'h0029,-16'h000b,16'h0021,16'h0059,16'h000f,16'h0016,16'h001a,-16'h003c,-16'h0010,-16'h0021,-16'h0078,-16'h001f,16'h004b,-16'h00a3,-16'h000e,16'h0068,16'h0001,16'h0001,16'h0000,-16'h000b,-16'h0022,16'h0014,-16'h0037,-16'h0076,16'h0064,16'h0004,16'h000a,16'h0019,-16'h0023,-16'h006b,16'h000b,16'h000c,16'h0037,16'h002f,-16'h0067,16'h0037,16'h0018,-16'h0008,16'h001f,16'h000f,16'h0000,-16'h002e,-16'h0008,16'h0024,-16'h0005,-16'h0052,16'h0023,-16'h006b,16'h002c,16'h00b6,-16'h0029,-16'h0074,16'h0036,16'h0014,16'h002e,16'h0023,16'h0052,-16'h003b,16'h0006,16'h0022,-16'h0033,16'h002c,-16'h004c,-16'h007e,-16'h0021,-16'h0019,16'h001b,16'h0063,16'h004c,16'h001f,16'h002b,-16'h0027,-16'h0028,-16'h0022,-16'h0067,16'h0016,16'h005a,-16'h00d0,-16'h0010,16'h0091,16'h0005,-16'h0007,16'h000b,-16'h0046,-16'h001f,16'h000f,-16'h0053,-16'h009e,16'h005f,-16'h0008,16'h001a,16'h0007,-16'h0051,-16'h007a,16'h0012,16'h0020,16'h0014,16'h0030,-16'h0083,-16'h0020,16'h0019,16'h0010,16'h001a,16'h000b,-16'h0017,-16'h000f,16'h0008,16'h001c,16'h0028,-16'h004d,16'h002a,-16'h0044,16'h0020,16'h00bf,-16'h0019,-16'h0073,16'h0051,16'h002a,16'h0038,16'h0011,16'h0039,-16'h0060,16'h000d,-16'h0004,-16'h0042,16'h001a,-16'h0080,-16'h0047,-16'h0029,16'h000d,16'h0011,16'h0047,16'h0045,16'h0006,16'h002e,-16'h0021,-16'h0026,-16'h0035,-16'h0074,16'h000d,16'h005c,-16'h010e,-16'h001d,16'h009d,16'h000c,-16'h000a,16'h0027,-16'h0038,-16'h001e,-16'h0003,-16'h0053,-16'h0078,16'h0034,16'h0014,16'h0021,-16'h0008,-16'h0041,-16'h0055,16'h0021,16'h002a,16'h0023,16'h0037,-16'h0069,-16'h008c,16'h0032,16'h0003,16'h003d,16'h0019,-16'h000e,16'h0006,-16'h0021,16'h003e,16'h001c,-16'h0051,16'h002e,-16'h0028,16'h0021,16'h00a2,-16'h001b,-16'h00bd,16'h006f,16'h004c,-16'h0003,16'h0021,16'h001c,-16'h0056,-16'h0013,16'h0020,-16'h007d,-16'h000e,-16'h0095,16'h0009,-16'h000c,16'h0021,16'h0035,16'h0023,16'h0044,16'h0023,16'h002a,16'h000c,-16'h0014,-16'h0023,-16'h005c,16'h0010,16'h006e,-16'h0114,16'h000c,16'h0091,16'h0021,-16'h0011,16'h0010,-16'h002a,-16'h0013,16'h0000,-16'h0051,-16'h0066,16'h001d,16'h0010,16'h0004,16'h000a,-16'h004d,-16'h0045,16'h002b,16'h0020,16'h002b,16'h005a,-16'h0076,-16'h00db,16'h004a,-16'h000d,16'h001f,16'h0048,-16'h001b,16'h0038,-16'h002b,16'h005f,16'h0013,-16'h006e,16'h0021,16'h0006,-16'h0021,16'h0097,-16'h001e,-16'h00ab,16'h005d,16'h0022,16'h0000,16'h001e,16'h0016,-16'h0072,-16'h001f,-16'h000f,-16'h00a4,16'h0007,-16'h0080,-16'h0016,-16'h0011,16'h0003,16'h000d,16'h000d,16'h0061,16'h0008,16'h0042,16'h0018,-16'h001f,-16'h0015,-16'h0054,-16'h0003,16'h0043,-16'h00e1,16'h000e,16'h0086,16'h0021,-16'h0010,-16'h0015,-16'h0027,-16'h0008,-16'h0027,-16'h003b,-16'h002e,-16'h0001,-16'h0015,-16'h0004,-16'h0001,-16'h0047,-16'h003b,16'h0004,16'h0014,-16'h0006,16'h006b,-16'h0067,-16'h00fe,16'h004b,-16'h002c,16'h000d,16'h004c,-16'h0019,16'h0017,-16'h001a,16'h0079,16'h0012,-16'h004f,-16'h0024,16'h0020,-16'h0031,16'h009a,-16'h0018,-16'h00d1,16'h004e,16'h000f,16'h0009,16'h001f,16'h0018,-16'h0095,-16'h003a,16'h0007,-16'h007a,16'h0005,-16'h004f,16'h0013,-16'h000a,16'h001f,16'h003a,16'h0049,16'h006b,-16'h0010,16'h0032,16'h0020,-16'h0013,16'h001c,-16'h003b,16'h001d,16'h0033,-16'h00d4,-16'h000c,16'h0087,16'h0003,-16'h0041,-16'h0016,-16'h0003,16'h0016,16'h0012,-16'h0040,16'h000f,-16'h002c,16'h000e,-16'h002e,16'h003e,-16'h0063,-16'h0013,16'h0024,16'h001f,-16'h0005,16'h0051,-16'h0061,-16'h011a,16'h003f,16'h0000,16'h0032,16'h003d,-16'h002a,16'h0012,-16'h003f,16'h006e,16'h0004,-16'h0072,16'h0000,16'h0035,-16'h0027,16'h008d,-16'h0001,-16'h00ed,16'h005f,-16'h0003,16'h001a,16'h002e,-16'h0007,-16'h00c6,-16'h0075,16'h0004,-16'h0063,-16'h000e,-16'h0035,-16'h000e,16'h001d,16'h002f,16'h0038,16'h0011,16'h0067,-16'h0023,16'h0056,16'h0016,-16'h0042,-16'h0007,-16'h0031,-16'h000b,16'h001c,-16'h00ab,-16'h0018,16'h008d,16'h0000,-16'h0042,-16'h0009,-16'h0008,16'h0065,-16'h0005,-16'h0021,16'h0033,-16'h0044,16'h0015,-16'h005f,16'h0025,-16'h0043,-16'h001b,16'h0007,-16'h0009,16'h0002,16'h003a,-16'h006d,-16'h0111,16'h0030,-16'h0003,16'h0019,16'h0051,-16'h0027,-16'h0011,-16'h0010,16'h005c,16'h000b,-16'h0076,-16'h0024,16'h004e,-16'h002c,16'h006d,16'h0019,-16'h00e9,16'h0056,16'h000b,16'h0000,16'h0007,-16'h0033,-16'h00e7,-16'h00b4,16'h001a,-16'h0097,-16'h0011,16'h0000,-16'h0002,16'h0014,16'h0017,16'h001c,16'h0003,16'h0019,-16'h002d,16'h004b,-16'h000b,-16'h0013,16'h0002,-16'h003b,16'h0007,16'h0040,-16'h00a4,-16'h005b,16'h0075,-16'h0008,-16'h005d,16'h0018,16'h0011,16'h0080,16'h0021,-16'h0007,16'h0030,-16'h0026,-16'h0001,-16'h0058,16'h003d,-16'h004a,-16'h002a,16'h0000,-16'h0004,16'h0015,16'h0014,-16'h0071,-16'h00f1,16'h0032,-16'h0001,16'h001e,16'h002f,-16'h0023,-16'h0021,-16'h0038,16'h0065,16'h0013,-16'h0055,-16'h0010,16'h005e,-16'h0003,16'h0086,16'h001a,-16'h00b0,16'h0071,16'h0016,16'h0011,16'h0027,-16'h002e,-16'h0114,-16'h00d6,16'h0012,-16'h0089,-16'h0022,-16'h0023,-16'h000f,16'h0033,-16'h0006,16'h0022,-16'h0012,-16'h0048,-16'h002c,16'h005c,-16'h0014,-16'h0017,16'h000e,-16'h0027,16'h0000,16'h0030,-16'h0072,-16'h00a5,16'h0078,-16'h0015,-16'h0046,16'h0014,16'h000b,16'h0092,16'h0024,-16'h0009,16'h0042,-16'h0044,16'h001e,-16'h0017,16'h0038,-16'h0041,-16'h000c,16'h0028,-16'h0006,16'h0015,16'h000a,-16'h0079,-16'h00a7,16'h0048,-16'h0003,16'h003f,16'h001d,-16'h0025,-16'h0031,16'h0004,16'h0048,16'h0007,-16'h002e,-16'h0022,16'h006d,16'h000b,16'h006e,16'h0035,-16'h00e1,16'h0061,16'h003a,16'h001e,16'h0006,-16'h003e,-16'h0120,-16'h0107,16'h0013,-16'h009b,-16'h0046,-16'h000c,-16'h003a,16'h0028,16'h0019,16'h0020,-16'h001d,-16'h0042,-16'h0020,16'h006a,-16'h0030,-16'h0024,16'h0011,-16'h0038,16'h001f,16'h0028,-16'h0046,-16'h00cd,16'h0064,-16'h001f,-16'h003a,16'h0016,-16'h0013,16'h0089,16'h002c,-16'h0019,16'h0062,-16'h0019,16'h001f,16'h000f,16'h0042,-16'h0014,-16'h000f,-16'h000d,16'h0009,16'h0006,16'h0016,-16'h005b,-16'h0090,16'h002f,16'h0017,16'h0020,16'h001a,-16'h0045,-16'h005e,16'h0012,16'h004d,-16'h000b,-16'h0014,-16'h0013,16'h005b,16'h0017,16'h0072,16'h0027,-16'h00d3,16'h004c,16'h0014,16'h0031,16'h002a,-16'h0069,-16'h013a,-16'h00c4,16'h000a,-16'h00bf,-16'h003e,-16'h0017,-16'h001f,16'h0041,16'h003c,16'h000c,-16'h002f,-16'h0045,16'h0003,16'h0046,-16'h000c,-16'h0035,16'h001a,-16'h005d,-16'h000e,16'h0039,-16'h004f,-16'h00c3,16'h0063,-16'h0017,-16'h003d,16'h0019,16'h0008,16'h009a,16'h003f,-16'h0004,16'h0052,16'h0007,16'h002a,16'h004f,16'h003b,16'h000f,-16'h0036,-16'h0011,16'h0000,16'h0000,-16'h0015,-16'h0043,-16'h005d,-16'h0008,16'h0011,16'h0056,16'h0016,-16'h001f,-16'h0076,16'h0028,16'h0070,-16'h0009,-16'h0015,-16'h0002,16'h0042,16'h003a,16'h004e,16'h0032,-16'h00c1,16'h0058,16'h0030,16'h0038,16'h0042,-16'h0087,-16'h0113,-16'h00a9,16'h0005,-16'h00bd,-16'h005f,-16'h0011,-16'h002d,16'h002d,16'h000d,16'h0018,-16'h001b,-16'h003a,16'h0008,16'h0029,-16'h0002,-16'h003a,16'h002b,-16'h004c,-16'h000b,16'h0033,-16'h0049,-16'h009b,16'h0054,-16'h0015,-16'h005d,-16'h0001,16'h000b,16'h00ac,16'h0003,-16'h001b,16'h0053,16'h0012,16'h002f,16'h0044,-16'h000a,16'h000b,-16'h004d,16'h000e,-16'h000e,16'h0023,-16'h006f,-16'h0012,-16'h001a,16'h0026,16'h000c,16'h0022,-16'h0004,16'h0000,-16'h0053,16'h0037,16'h005d,-16'h000a,-16'h0041,16'h000b,16'h002e,16'h0045,16'h0089,16'h001c,-16'h0088,16'h006c,16'h0033,16'h0021,16'h0037,-16'h0096,-16'h011b,-16'h0090,16'h0010,-16'h007a,-16'h006d,-16'h0012,-16'h0018,16'h0027,16'h000c,16'h0018,16'h000e,-16'h002f,16'h0021,16'h002d,16'h0007,-16'h0036,16'h003b,-16'h003d,-16'h001b,16'h0018,-16'h0031,-16'h006c,16'h0022,16'h0009,-16'h0060,16'h0020,16'h001d,16'h00c5,16'h0001,-16'h0033,16'h002e,16'h001a,16'h0030,16'h0035,-16'h0018,-16'h0010,-16'h004b,16'h0003,16'h000a,16'h0014,-16'h00e7,16'h0012,-16'h000a,-16'h000f,16'h0012,16'h0035,16'h0023,-16'h000d,16'h0001,16'h0028,16'h0058,-16'h000a,-16'h0058,16'h0036,16'h0025,16'h005d,16'h0054,-16'h0024,-16'h008e,16'h008f,16'h003c,16'h0029,16'h0056,-16'h00c4,-16'h00d7,-16'h0046,16'h0010,-16'h007b,-16'h005a,-16'h0010,-16'h0010,16'h0030,16'h0010,16'h001c,16'h0010,16'h000c,16'h002a,16'h0011,16'h0040,-16'h0032,16'h002e,-16'h004f,-16'h000a,16'h0023,-16'h001e,-16'h004e,16'h0020,-16'h000b,-16'h004c,16'h0029,16'h001c,16'h00e5,16'h000a,-16'h001c,16'h000a,16'h001c,16'h001c,16'h001d,-16'h0027,-16'h0008,-16'h0041,16'h0035,-16'h0009,16'h0023,-16'h012e,16'h0032,-16'h0010,16'h0008,16'h0002,16'h002a,-16'h0005,-16'h0013,16'h001d,16'h0038,16'h0070,-16'h000e,-16'h005c,16'h003b,16'h0027,16'h0019,16'h0061,-16'h0029,-16'h00af,16'h0078,16'h0031,16'h002a,16'h0040,-16'h00e6,-16'h00a0,-16'h0007,-16'h0019,-16'h0088,-16'h006f,16'h0002,16'h0012,16'h0006,16'h001a,16'h0009,16'h0025,16'h0024,16'h0034,-16'h0021,16'h0042,-16'h002b,16'h0015,-16'h002b,16'h002d,-16'h001e,-16'h0008,-16'h0035,16'h002f,-16'h0012,-16'h004c,16'h0030,16'h000f,16'h00ae,16'h001b,-16'h000d,16'h000d,16'h001a,16'h0028,16'h0039,-16'h0066,16'h000e,-16'h0056,16'h0044,16'h0014,16'h001b,-16'h012d,16'h0074,-16'h000a,16'h0000,-16'h0022,16'h0005,16'h000b,16'h0001,16'h0028,16'h0030,16'h0030,-16'h0072,-16'h007d,16'h002d,16'h000b,16'h0005,16'h0025,-16'h002c,-16'h00a7,16'h0092,16'h0023,16'h0024,16'h0037,-16'h00ed,-16'h0042,-16'h0012,-16'h0010,-16'h0061,-16'h0064,16'h0042,-16'h000d,16'h0034,16'h0012,16'h0005,16'h0040,16'h0064,16'h0016,-16'h0016,16'h005b,-16'h002e,16'h003b,-16'h0043,16'h001f,-16'h0018,16'h0007,-16'h0039,16'h0027,-16'h001c,-16'h0078,16'h0006,-16'h0004,16'h0052,-16'h0005,-16'h000c,16'h000d,16'h0017,16'h0043,16'h0040,-16'h00c6,16'h0018,16'h0002,-16'h0001,16'h0000,16'h0012,-16'h00e8,16'h0067,16'h0013,-16'h000f,-16'h0022,16'h0022,16'h002a,16'h002d,16'h0039,16'h0006,-16'h0005,-16'h0078,-16'h004f,16'h0007,-16'h0005,-16'h0013,16'h000d,16'h0012,-16'h00c5,16'h0093,16'h0022,16'h0045,16'h002b,-16'h00c8,-16'h001a,16'h0009,-16'h0019,-16'h0057,-16'h008a,16'h005c,-16'h0009,16'h001d,16'h0041,-16'h0005,16'h0051,16'h0057,16'h002e,-16'h0006,16'h007d,16'h0002,16'h0051,-16'h003e,16'h0015,-16'h0025,16'h004a,-16'h002e,16'h001e,-16'h0032,-16'h006d,16'h0016,16'h000e,16'h0014,16'h0007,-16'h000b,-16'h0031,16'h001a,16'h005f,16'h001c,-16'h0109,16'h0040,16'h0034,16'h0015,-16'h0016,16'h0013,-16'h0091,16'h0085,16'h0024,-16'h001f,-16'h001b,-16'h0013,16'h000b,16'h0002,16'h002a,16'h000b,-16'h0021,-16'h007d,-16'h0033,16'h0019,16'h0002,-16'h0033,16'h0016,16'h003e,-16'h00bd,16'h00af,16'h0023,16'h0022,16'h0030,-16'h00ab,-16'h0002,16'h0037,-16'h0037,-16'h005f,-16'h0082,16'h0052,-16'h0037,16'h0036,16'h005b,16'h0014,16'h0046,16'h004e,16'h0013,16'h0007,16'h007b,-16'h0014,16'h0064,-16'h0042,16'h0021,-16'h001e,16'h0040,-16'h003c,16'h0022,-16'h0037,-16'h0054,16'h0015,-16'h0026,-16'h0017,16'h003a,16'h000d,-16'h004f,16'h0016,16'h004e,16'h0005,-16'h00ac,16'h0030,16'h003a,-16'h0001,-16'h001d,16'h0017,-16'h006d,16'h0079,16'h0016,-16'h002f,-16'h0048,-16'h0019,16'h0020,16'h0003,16'h0006,-16'h000b,-16'h006d,-16'h009e,-16'h0036,-16'h001c,16'h0019,-16'h0056,16'h0022,16'h006d,-16'h00c2,16'h00a1,16'h0037,16'h0031,16'h0022,-16'h0076,16'h000b,16'h004e,-16'h003e,-16'h0068,-16'h0067,16'h006f,-16'h0045,16'h0027,16'h005d,-16'h001e,16'h004b,16'h0044,16'h0015,16'h0006,16'h0057,16'h0021,16'h006a,-16'h004d,16'h0030,-16'h0008,16'h001f,-16'h0035,16'h0038,-16'h0026,-16'h0047,-16'h0008,-16'h000c,-16'h0050,16'h0017,16'h0023,-16'h0084,16'h002d,16'h004e,-16'h003a,-16'h0088,16'h0058,16'h0045,16'h0008,-16'h004a,16'h002b,-16'h0020,16'h0080,16'h0029,-16'h002b,-16'h006f,-16'h0015,16'h002d,16'h0011,-16'h0029,-16'h0008,-16'h0052,-16'h0052,-16'h0051,-16'h0050,16'h002e,-16'h0068,16'h004f,16'h0064,-16'h00a5,16'h008c,16'h006d,16'h0002,16'h0039,-16'h0060,-16'h0011,16'h005e,-16'h003e,-16'h0058,-16'h0070,16'h0056,-16'h001e,16'h000a,16'h0038,-16'h0022,16'h003d,16'h0024,16'h0005,16'h002c,16'h0048,16'h0057,16'h003e,-16'h004d,16'h0003,16'h0029,16'h0025,-16'h001b,16'h001f,-16'h0004,-16'h0041,-16'h0008,-16'h0004,-16'h0042,16'h0027,16'h0033,-16'h00c3,16'h002c,16'h003e,-16'h0024,-16'h001e,16'h0061,16'h0018,16'h0016,-16'h003c,16'h000c,-16'h001e,16'h0085,16'h003a,-16'h000c,-16'h0077,-16'h0026,16'h0049,16'h0016,-16'h0034,16'h001a,-16'h0030,-16'h0044,-16'h0043,-16'h004c,16'h005f,-16'h0049,16'h0075,16'h006a,-16'h005f,16'h006a,16'h0059,16'h001f,16'h0030,-16'h0021,16'h000f,16'h004e,-16'h003f,-16'h004b,-16'h004a,16'h003e,-16'h0022,16'h0000,16'h0004,-16'h001b,16'h0028,16'h001b,-16'h0012,16'h003e,16'h0018,16'h0043,16'h002a,-16'h004f,-16'h001b,16'h0021,16'h001b,-16'h0011,16'h0014,-16'h000d,-16'h0025,16'h0026,-16'h0010,-16'h0027,16'h000d,16'h0022,-16'h00af,16'h001a,16'h0042,-16'h001e,16'h0017,16'h004d,16'h001a,16'h000f,-16'h0031,16'h0026,-16'h0002,16'h0056,16'h000c,-16'h0028,-16'h004c,16'h0009,16'h000a,-16'h000b,-16'h0036,16'h0028,-16'h0028,-16'h0046,-16'h0025,-16'h002e,16'h004a,-16'h0031,16'h0083,16'h003f,-16'h003d,16'h005f,16'h0079,16'h001d,16'h0068,-16'h002b,-16'h0001,16'h0052,16'h0009,-16'h0041,-16'h003a,16'h003c,16'h0000,-16'h000c,16'h000d,-16'h0004,16'h002b,16'h0022,16'h000f,16'h0003,16'h000d,16'h004e,16'h0024,-16'h0034,16'h0005,16'h0065,16'h000c,16'h0009,16'h0038,-16'h0005,-16'h001d,16'h0044,-16'h0008,-16'h000b,16'h0015,16'h0047,-16'h00af,-16'h0013,16'h0017,-16'h0012,16'h0003,16'h0068,16'h0011,16'h0014,-16'h0032,16'h0033,16'h000d,16'h0061,16'h0029,-16'h0022,-16'h0051,16'h0015,16'h001c,-16'h0007,-16'h0026,16'h002a,-16'h0029,-16'h000d,-16'h0035,-16'h001d,16'h002b,-16'h0022,16'h0072,16'h0009,-16'h0013,16'h0037,16'h0090,-16'h0007,16'h0073,-16'h000d,16'h0026,16'h0019,-16'h000e,-16'h0020,16'h001a,16'h0071,-16'h002a,-16'h0003,16'h0004,-16'h0005,16'h0007,16'h0014,16'h001f,-16'h0014,-16'h0011,16'h0046,16'h0028,-16'h001f,16'h0026,16'h0056,-16'h000e,16'h0012,16'h0057,16'h0011,16'h0005,16'h0047,-16'h0003,-16'h000a,-16'h0019,16'h0037,-16'h009b,-16'h0020,16'h0024,-16'h000c,16'h0014,16'h004c,-16'h000e,16'h0015,-16'h002d,16'h0044,-16'h0005,16'h002e,16'h0017,-16'h0043,-16'h003b,16'h0005,16'h0017,16'h0004,-16'h0012,16'h0018,-16'h0007,-16'h0021,-16'h0042,-16'h0022,16'h005f,-16'h001c,16'h0052,-16'h002d,-16'h001f,16'h0048,16'h007f,-16'h001f,16'h007b,-16'h0004,16'h0058,16'h000c,-16'h000a,-16'h001e,16'h0046,16'h006e,-16'h003b,16'h0008,16'h0028,16'h0011,16'h0017,-16'h0005,-16'h0010,-16'h0022,-16'h001f,16'h003d,16'h0022,16'h0002,16'h0015,16'h000d,-16'h0020,-16'h0029,16'h0019,16'h0012,-16'h0013,16'h000f,16'h0055,-16'h004c,16'h000f,-16'h0007,-16'h000a,16'h004b,-16'h000f,-16'h0081,-16'h000f,16'h0065,-16'h0011,16'h0025,-16'h0012,16'h003d,-16'h0001,-16'h0014,16'h0021,16'h0019,-16'h0042,16'h0016,-16'h000c,16'h001c,-16'h0026,-16'h0004,-16'h002a,-16'h0057,-16'h0033,-16'h0025,-16'h001d,-16'h0021,16'h006f,-16'h0022,-16'h0017,16'h0035,-16'h0010,16'h0060,16'h0027,16'h0027,-16'h0017,-16'h0033,16'h004d,-16'h0001,16'h0020,-16'h0018,-16'h0004,-16'h0016,-16'h003f,16'h0007,16'h0054,-16'h007a,16'h0039,16'h0022,16'h0038,-16'h0002,-16'h0020,-16'h003f,-16'h002f,-16'h0019,-16'h0020,-16'h001f,16'h003a,16'h0031,16'h000e,-16'h001c,16'h000f,-16'h0079,16'h0010,16'h0002,-16'h000c,16'h0049,16'h0002,-16'h0089,16'h001d,16'h004c,16'h000b,16'h000f,16'h001a,16'h001d,-16'h0003,-16'h002e,16'h0068,16'h0011,-16'h0050,16'h0030,16'h0011,16'h0007,-16'h0001,16'h0012,-16'h0025,-16'h0028,-16'h000d,-16'h0005,-16'h0018,16'h001a,16'h0069,16'h0027,-16'h0040,16'h0033,-16'h003c,16'h005b,16'h002a,16'h0033,-16'h0017,-16'h0013,16'h002c,16'h000a,-16'h0007,-16'h0029,-16'h0029,-16'h0029,16'h0002,16'h0004,16'h004d,-16'h0061,16'h000b,-16'h000d,16'h0002,-16'h0013,-16'h0034,-16'h004d,-16'h0051,16'h000e,-16'h002b,16'h0001,16'h0049,16'h0024,-16'h000d,-16'h0003,16'h0010,-16'h009a,16'h001a,16'h001e,-16'h001f,16'h0045,16'h000e,-16'h0070,16'h002b,16'h0052,-16'h0005,16'h0019,-16'h0004,16'h0024,-16'h0007,-16'h0030,16'h00ab,16'h000c,-16'h0047,16'h0023,16'h0008,16'h0019,-16'h000d,16'h0007,-16'h002f,-16'h0017,-16'h0014,-16'h0007,-16'h003a,-16'h0001,16'h009b,16'h000e,-16'h004a,16'h0051,-16'h002e,16'h004f,16'h0022,16'h0046,-16'h0013,-16'h0008,16'h002e,-16'h0030,16'h0005,-16'h004b,-16'h006a,-16'h002d,-16'h001b,-16'h0012,16'h0039,-16'h0023,16'h002e,-16'h000d,-16'h001b,-16'h0012,-16'h004c,-16'h005a,-16'h0075,16'h0023,-16'h0064,16'h0015,16'h004a,16'h000b,-16'h002d,-16'h0029,16'h0017,-16'h007e,16'h000e,16'h000e,-16'h0059,16'h005b,16'h0004,-16'h003a,16'h0042,16'h002e,-16'h0012,-16'h0005,16'h0006,16'h0035,16'h0009,-16'h0055,16'h008f,16'h002c,-16'h002d,16'h0020,16'h0003,16'h0016,16'h0003,16'h0025,-16'h000e,-16'h0017,16'h0004,16'h0031,-16'h0061,16'h0019,16'h00b9,16'h0005,-16'h006c,16'h003e,-16'h0024,16'h0055,16'h001b,16'h004d,-16'h001f,16'h0020,16'h0048,-16'h0036,16'h001e,-16'h004a,-16'h0090,-16'h004a,-16'h000f,-16'h0033,16'h005e,-16'h0003,16'h0018,16'h000a,-16'h004c,16'h0007,-16'h000d,-16'h004a,-16'h0028,16'h0039,-16'h006b,16'h0027,16'h0053,-16'h0020,-16'h0020,-16'h0010,16'h0012,-16'h0060,16'h0031,16'h000c,-16'h006b,16'h0046,16'h0005,16'h0028,16'h003a,-16'h001b,16'h0002,-16'h000c,-16'h001f,16'h002b,-16'h001a,-16'h006d,16'h0081,16'h0016,-16'h000b,16'h001c,-16'h0020,16'h000e,-16'h001e,16'h0031,16'h0014,16'h0014,-16'h0045,16'h0033,-16'h0056,16'h0009,16'h009b,-16'h0011,-16'h0066,16'h0031,16'h0005,16'h0039,16'h003c,16'h004c,-16'h0022,16'h0012,16'h0007,-16'h0043,16'h0058,-16'h008b,-16'h0096,-16'h0034,-16'h0017,-16'h0024,16'h004e,16'h003b,16'h0038,16'h0013,-16'h0056,16'h0002,-16'h003a,-16'h0044,-16'h0009,16'h005d,-16'h00b3,16'h0007,16'h0061,-16'h0024,16'h0009,16'h0015,-16'h0011,-16'h0029,16'h0032,-16'h0004,-16'h008f,16'h0061,-16'h0010,16'h001f,16'h0016,-16'h0069,-16'h001c,16'h001d,16'h0005,16'h004a,16'h001e,-16'h0043,16'h002b,16'h0005,-16'h0006,16'h0036,-16'h0010,16'h0018,-16'h000a,16'h0035,16'h0034,16'h001b,-16'h004b,16'h0021,-16'h0068,16'h0009,16'h00a2,-16'h0021,-16'h0069,16'h004b,16'h0024,16'h0041,16'h002c,16'h004e,-16'h002d,16'h0023,-16'h0007,-16'h0051,16'h0048,-16'h0092,-16'h0042,-16'h004c,16'h000c,-16'h0016,16'h0042,16'h003a,16'h0038,16'h0034,-16'h0040,16'h0012,-16'h0030,-16'h004e,16'h0009,16'h0061,-16'h00b6,16'h0014,16'h0077,-16'h0007,-16'h001c,-16'h0009,-16'h0035,-16'h0026,16'h0011,-16'h002f,-16'h009e,16'h0051,16'h0012,16'h0044,-16'h0002,-16'h0072,-16'h0010,16'h0013,-16'h0005,16'h0014,16'h0029,-16'h0053,-16'h0056,16'h001f,16'h0002,16'h0058,16'h0003,-16'h0006,16'h0012,-16'h0002,16'h0050,16'h0035,-16'h0063,16'h0034,-16'h0010,16'h0026,16'h0089,-16'h001f,-16'h006f,16'h0033,16'h003b,-16'h0006,16'h000c,16'h0037,-16'h003f,16'h0004,-16'h0022,-16'h0098,16'h002a,-16'h00ac,-16'h0005,-16'h004e,16'h000f,16'h0003,16'h004e,16'h002c,-16'h0002,16'h003a,16'h0006,16'h000b,-16'h0024,-16'h0023,16'h0004,16'h005c,-16'h009c,16'h0047,16'h007e,16'h0001,-16'h0006,-16'h0028,-16'h0043,-16'h002c,-16'h0016,-16'h0034,-16'h0087,16'h004c,-16'h0007,16'h0035,16'h000f,-16'h006b,-16'h002d,16'h000b,16'h0013,16'h0019,16'h0023,-16'h0045,-16'h00c0,16'h000c,-16'h0005,16'h0039,16'h0011,16'h0008,16'h0019,16'h0017,16'h0022,16'h002a,-16'h0067,16'h0005,16'h0009,16'h000f,16'h0074,-16'h0013,-16'h008b,16'h0055,16'h000d,16'h0006,16'h000c,16'h0046,-16'h0051,16'h0000,-16'h0001,-16'h00ba,16'h0005,-16'h0089,16'h0005,-16'h003c,16'h004d,-16'h0008,16'h004e,16'h0052,16'h0005,16'h003c,16'h0005,16'h0008,-16'h0011,-16'h001d,16'h0011,16'h004c,-16'h0075,16'h003f,16'h0097,16'h000e,-16'h0006,-16'h0008,-16'h0032,16'h0013,-16'h001f,-16'h0044,-16'h0076,16'h0023,-16'h0015,16'h002f,16'h0007,-16'h0024,-16'h0012,16'h000c,16'h0003,16'h0007,16'h002c,-16'h0058,-16'h00e9,16'h0041,-16'h001a,16'h0030,16'h0017,-16'h0027,16'h000a,-16'h0005,16'h006e,-16'h0006,-16'h006c,16'h0004,16'h001d,-16'h0032,16'h0071,-16'h003c,-16'h0082,16'h004d,16'h0024,-16'h0003,16'h0027,16'h0019,-16'h0077,-16'h0033,-16'h001e,-16'h00a5,-16'h0021,-16'h006b,16'h0005,-16'h001c,16'h003b,16'h0020,16'h0032,16'h003d,16'h0007,16'h0044,16'h0021,16'h0017,16'h0005,-16'h001a,16'h0018,16'h004e,-16'h0056,16'h0020,16'h00a4,16'h0000,-16'h0003,-16'h0017,-16'h0009,16'h000b,-16'h0013,-16'h0040,-16'h0040,-16'h000a,-16'h000f,-16'h0013,16'h0000,-16'h003c,-16'h0002,-16'h000f,-16'h0009,16'h0013,16'h0030,-16'h0035,-16'h012b,16'h0020,-16'h000c,16'h0023,16'h0028,-16'h0027,16'h002d,-16'h001f,16'h0053,16'h000e,-16'h005e,16'h0000,16'h0049,-16'h0033,16'h007b,-16'h0013,-16'h009e,16'h0043,16'h0001,-16'h001c,16'h0041,-16'h000a,-16'h0076,-16'h0053,-16'h0030,-16'h007b,-16'h001a,-16'h0026,-16'h0010,-16'h0019,16'h001c,16'h000b,16'h001b,16'h0038,-16'h0023,16'h0015,16'h0007,16'h000d,16'h0022,-16'h0028,16'h0016,16'h0043,-16'h0035,16'h0007,16'h0095,-16'h0003,-16'h0002,-16'h001a,-16'h0022,16'h003d,16'h000b,-16'h0034,-16'h0024,-16'h0027,-16'h0012,-16'h001d,16'h0013,-16'h0046,16'h000a,16'h000c,16'h0003,16'h0000,16'h0029,-16'h004f,-16'h0107,16'h0013,-16'h0001,16'h0018,16'h003b,-16'h0001,16'h0013,-16'h003b,16'h006b,-16'h0005,-16'h003f,-16'h0012,16'h0056,-16'h0039,16'h008d,16'h000b,-16'h009e,16'h005f,-16'h000d,16'h0003,16'h002b,-16'h001e,-16'h009c,-16'h0072,-16'h0018,-16'h0082,-16'h002d,-16'h0006,-16'h0009,-16'h0016,16'h0026,-16'h0001,-16'h0008,16'h0006,-16'h0014,16'h0035,-16'h0029,-16'h0002,16'h0009,-16'h0011,-16'h0034,16'h0006,-16'h0048,-16'h0019,16'h0084,-16'h001b,16'h0017,-16'h0016,16'h0001,16'h003c,16'h000e,-16'h0037,-16'h0016,-16'h002f,-16'h0004,-16'h0041,16'h001b,-16'h0050,16'h0003,-16'h001c,-16'h0020,-16'h000e,16'h0043,-16'h0037,-16'h00d4,16'h001e,16'h000a,16'h001b,16'h0054,-16'h0009,16'h000f,-16'h0028,16'h004a,-16'h0007,-16'h0048,-16'h0018,16'h0060,-16'h0004,16'h008d,16'h0007,-16'h009f,16'h0053,-16'h0007,16'h0012,16'h001d,-16'h0022,-16'h00cd,-16'h00a3,-16'h0018,-16'h0087,-16'h0038,16'h0007,-16'h0008,16'h0009,16'h001d,16'h0010,-16'h0007,-16'h0031,-16'h0037,16'h0030,-16'h002f,-16'h0009,16'h0031,-16'h002a,-16'h0007,16'h001b,-16'h0036,-16'h0040,16'h0057,-16'h0001,16'h001a,-16'h0008,16'h0016,16'h0077,16'h0021,-16'h0015,-16'h001e,-16'h0022,16'h0011,16'h0000,16'h0025,-16'h002f,-16'h0004,-16'h0017,-16'h0022,16'h0009,16'h004d,-16'h0049,-16'h0098,16'h000b,-16'h0005,16'h0009,16'h002a,-16'h0017,-16'h000e,-16'h003d,16'h003d,16'h0005,-16'h002b,-16'h0008,16'h005c,-16'h0006,16'h0073,16'h000f,-16'h00a2,16'h0041,-16'h000c,16'h0009,16'h0020,-16'h001b,-16'h0122,-16'h00ed,-16'h0027,-16'h0098,-16'h0034,-16'h0013,-16'h0008,16'h0014,16'h0023,16'h000c,-16'h001c,-16'h0083,-16'h0019,16'h0023,-16'h001c,16'h0008,-16'h000a,-16'h0022,-16'h000e,16'h0036,16'h0004,-16'h005f,16'h0065,16'h0010,16'h000d,-16'h0009,16'h001d,16'h008a,16'h0018,-16'h000a,16'h001e,-16'h002c,16'h001b,16'h0027,16'h0039,-16'h001a,-16'h0007,-16'h0030,-16'h0013,16'h000f,16'h0046,-16'h005c,-16'h004a,16'h0001,16'h0024,16'h001a,16'h003a,-16'h0028,-16'h000f,-16'h0009,16'h0030,16'h000e,-16'h0020,-16'h0007,16'h0056,16'h0000,16'h007e,16'h002a,-16'h00a7,16'h005d,16'h0017,-16'h000c,16'h000a,-16'h001d,-16'h0109,-16'h00de,-16'h0009,-16'h00a4,-16'h0052,-16'h0003,-16'h0023,16'h0018,16'h002e,16'h003e,-16'h001b,-16'h0075,-16'h0008,16'h0051,-16'h001e,-16'h0004,-16'h0009,-16'h0038,-16'h0001,16'h000c,16'h0009,-16'h0098,16'h0058,16'h0015,16'h0019,16'h000e,16'h002f,16'h0071,16'h0011,-16'h0003,16'h0039,-16'h0027,16'h0002,16'h0064,16'h0014,-16'h0003,-16'h0002,-16'h002a,16'h0007,16'h0023,16'h0044,-16'h001c,-16'h0019,-16'h000a,16'h000c,16'h002a,16'h000f,-16'h001f,-16'h0037,16'h0002,16'h002b,16'h0003,-16'h0025,-16'h000e,16'h0025,16'h000b,16'h008c,16'h003c,-16'h008e,16'h0056,16'h002d,-16'h0013,16'h0031,-16'h0012,-16'h00ef,-16'h00e0,-16'h0002,-16'h00a3,-16'h0082,-16'h001a,-16'h000f,16'h002a,16'h0024,16'h0034,-16'h0028,-16'h004d,16'h0005,16'h002c,-16'h000d,16'h0000,16'h0009,-16'h0038,-16'h001d,-16'h0002,16'h0025,-16'h006d,16'h0066,-16'h0019,-16'h0012,-16'h000e,16'h001d,16'h0080,16'h000a,16'h000a,16'h0049,-16'h0033,16'h0027,16'h0055,16'h0012,16'h000a,-16'h0017,-16'h0035,-16'h0009,16'h0013,16'h000b,-16'h0003,16'h0005,-16'h000a,16'h0014,16'h0016,-16'h000b,-16'h0011,-16'h004a,16'h000f,16'h0043,16'h0005,-16'h0017,16'h0006,16'h0002,16'h0032,16'h0077,16'h0048,-16'h0088,16'h0084,16'h0016,16'h000f,16'h003e,-16'h0033,-16'h00c9,-16'h00d8,16'h0021,-16'h009a,-16'h006c,-16'h0011,16'h0003,16'h0016,16'h0005,16'h0048,16'h000f,-16'h0018,16'h0013,16'h001f,16'h0019,-16'h0014,-16'h0003,-16'h003c,-16'h0019,-16'h000f,16'h0007,-16'h001d,16'h005f,-16'h000e,-16'h0038,16'h0003,16'h0005,16'h0093,-16'h0004,16'h0023,16'h004f,-16'h002c,16'h000a,16'h0024,16'h002a,-16'h0004,-16'h0026,-16'h0009,-16'h000f,-16'h0001,-16'h0018,16'h0010,16'h0034,-16'h001a,16'h0008,16'h0030,-16'h000b,16'h000e,-16'h003a,16'h0004,16'h004e,-16'h000c,-16'h0014,16'h0021,16'h0019,16'h0050,16'h008b,16'h0044,-16'h0067,16'h0079,16'h002c,-16'h0026,16'h001d,-16'h004d,-16'h00d6,-16'h00d4,16'h0016,-16'h007c,-16'h0059,16'h0003,16'h001a,16'h001f,-16'h0009,16'h005b,16'h001d,-16'h001c,16'h0022,-16'h0008,16'h001d,-16'h003a,16'h0032,-16'h000c,-16'h000c,16'h0006,-16'h0008,-16'h000d,16'h0046,16'h0010,-16'h007b,16'h000b,-16'h0002,16'h00a2,-16'h0011,16'h0010,16'h0047,16'h0007,-16'h002a,-16'h0007,16'h0048,-16'h0001,-16'h0024,-16'h0013,-16'h000e,16'h000a,-16'h00b0,16'h003a,16'h0031,-16'h004e,-16'h000d,16'h001f,-16'h002c,-16'h001b,-16'h0019,16'h000d,16'h0042,-16'h0004,-16'h0047,16'h0031,16'h0021,16'h0044,16'h007a,16'h0006,-16'h007d,16'h0077,16'h0030,-16'h001b,16'h0005,-16'h008f,-16'h00a3,-16'h009c,16'h0013,-16'h0062,-16'h0073,16'h0005,16'h0001,16'h000b,-16'h000f,16'h0044,16'h0030,16'h001f,16'h0017,16'h0001,16'h001b,-16'h0039,16'h0001,-16'h002b,-16'h0019,16'h0005,16'h0003,16'h0004,16'h0032,16'h000a,-16'h0047,16'h0000,16'h0015,16'h0090,-16'h0021,-16'h0008,16'h0021,16'h0007,-16'h0016,16'h0006,-16'h0018,16'h0019,-16'h003e,16'h0013,16'h0026,-16'h0007,-16'h012e,16'h004c,16'h001b,-16'h0039,-16'h001b,16'h0022,-16'h0023,-16'h000b,-16'h0002,16'h002a,16'h0039,-16'h0032,-16'h006a,16'h0026,16'h0010,16'h0049,16'h005a,-16'h0030,-16'h0060,16'h0081,16'h0021,16'h0002,16'h0016,-16'h00b7,-16'h005b,-16'h0052,16'h0035,-16'h0074,-16'h006f,16'h0004,16'h0013,16'h0038,-16'h0001,16'h004a,16'h0024,16'h0050,16'h0038,-16'h003f,16'h0036,-16'h0035,-16'h0003,-16'h002d,16'h0024,-16'h0001,16'h0002,-16'h0005,16'h0027,-16'h0002,-16'h004e,-16'h0007,-16'h0002,16'h005d,-16'h001b,-16'h0004,16'h0017,16'h001d,16'h000e,16'h0014,-16'h0041,16'h001c,-16'h0049,16'h0018,16'h0007,16'h001c,-16'h015d,16'h004a,-16'h0002,-16'h001f,-16'h0029,16'h0000,-16'h0021,-16'h000c,16'h0030,16'h0030,16'h000b,-16'h003d,-16'h0074,16'h001c,-16'h001b,16'h0026,16'h0039,-16'h0028,-16'h0052,16'h0090,16'h0023,16'h002d,16'h001d,-16'h00e0,-16'h001f,-16'h0047,16'h0016,-16'h0077,-16'h006d,16'h0000,16'h0018,16'h0031,-16'h0003,16'h003b,16'h003b,16'h004e,16'h000e,-16'h0031,16'h003a,-16'h001f,16'h000b,-16'h002b,16'h0031,-16'h0001,16'h0017,-16'h0019,16'h0024,-16'h0002,-16'h004b,-16'h0001,16'h0012,16'h0023,16'h0001,-16'h0009,-16'h0006,16'h0028,16'h0014,16'h001e,-16'h00bf,16'h002a,-16'h002f,-16'h000c,16'h0014,16'h0002,-16'h00f8,16'h004f,16'h0015,-16'h0017,-16'h0005,16'h0002,16'h0011,16'h001b,16'h005e,16'h0014,-16'h003d,-16'h0064,-16'h0045,-16'h000e,-16'h0030,16'h0007,16'h002a,16'h0000,-16'h0070,16'h00ae,16'h0007,16'h0034,16'h0002,-16'h00e8,16'h0013,-16'h0025,16'h0004,-16'h0080,-16'h006b,16'h003c,16'h000a,16'h0044,16'h0023,16'h0008,16'h001d,16'h0046,16'h0026,-16'h0033,16'h004c,-16'h0010,16'h0010,-16'h0017,16'h004e,16'h0001,16'h002a,-16'h0048,16'h0017,16'h000a,-16'h0030,-16'h0006,-16'h0009,-16'h0020,16'h0022,-16'h001c,-16'h0010,16'h0039,16'h0029,16'h0004,-16'h0155,16'h003b,-16'h0006,16'h0011,16'h0008,16'h0042,-16'h007c,16'h005e,16'h000f,16'h0017,-16'h0021,-16'h0014,16'h001a,16'h0013,16'h0034,-16'h0021,-16'h007a,-16'h0055,-16'h0028,-16'h0018,-16'h0015,-16'h003c,16'h0010,16'h0023,-16'h006f,16'h0089,16'h003d,16'h0037,-16'h001c,-16'h00dd,16'h0028,-16'h0009,16'h0016,-16'h0046,-16'h0082,16'h001c,16'h0003,16'h0024,16'h0046,-16'h0002,16'h003f,16'h0030,16'h003f,-16'h000f,16'h007a,16'h001d,16'h0002,-16'h0012,16'h004f,-16'h0010,16'h0053,-16'h0019,16'h0020,16'h002b,-16'h001a,16'h0001,-16'h0007,-16'h0049,16'h001c,-16'h001a,-16'h004d,16'h0054,16'h0030,-16'h002a,-16'h00fb,16'h002c,16'h0031,16'h001c,-16'h0016,16'h0057,-16'h0065,16'h0044,16'h001b,-16'h002b,-16'h002c,-16'h0001,16'h0032,16'h000e,16'h0016,-16'h003b,-16'h008b,-16'h0055,-16'h0026,-16'h001a,-16'h0001,-16'h0024,16'h001f,16'h008e,-16'h0058,16'h0087,16'h0027,16'h0038,-16'h0017,-16'h00a2,16'h002e,16'h0010,-16'h0026,-16'h005d,-16'h003e,16'h0038,-16'h0023,16'h0030,16'h0046,-16'h0011,16'h0040,16'h003f,16'h005b,16'h000a,16'h005a,16'h003d,16'h000a,-16'h0031,16'h0023,-16'h001f,16'h004f,16'h000b,16'h0030,16'h001e,-16'h0027,-16'h0007,-16'h000b,-16'h0066,16'h000a,-16'h0021,-16'h0092,16'h004e,16'h003e,-16'h0030,-16'h00a4,16'h0049,16'h0040,16'h000b,-16'h002e,16'h0018,-16'h002e,16'h003a,16'h002b,-16'h0034,-16'h004e,-16'h000a,16'h0037,16'h0006,16'h0008,-16'h0042,-16'h007e,-16'h0044,-16'h0043,16'h0002,16'h0003,-16'h002a,16'h0047,16'h0093,-16'h004c,16'h009c,16'h0043,16'h0039,-16'h0029,-16'h0065,16'h0045,16'h0033,-16'h0039,-16'h0067,-16'h0038,16'h0038,-16'h0015,16'h0029,16'h001c,-16'h0020,16'h0050,16'h0023,16'h0038,16'h003b,16'h0060,16'h0057,16'h0015,-16'h0046,16'h0030,16'h0018,16'h003c,16'h001f,16'h002c,16'h0017,-16'h001e,-16'h002d,-16'h001f,-16'h005e,-16'h0001,16'h001b,-16'h00d3,16'h0054,16'h003a,-16'h0036,-16'h0041,16'h002b,16'h0036,-16'h001e,-16'h0036,16'h000b,-16'h000a,16'h0044,16'h0019,-16'h004f,-16'h0054,-16'h0019,16'h001c,-16'h000d,16'h0010,-16'h001b,-16'h005d,-16'h004a,-16'h0057,-16'h0028,16'h000d,-16'h0051,16'h0076,16'h0091,-16'h0038,16'h008a,16'h0034,16'h0025,16'h0004,-16'h003a,16'h0044,16'h0041,-16'h0042,-16'h007b,-16'h0029,16'h004f,-16'h002e,16'h0005,16'h0000,-16'h0043,16'h0012,16'h001c,16'h0013,16'h006d,16'h0024,16'h0075,16'h0008,-16'h003c,16'h0022,16'h0023,16'h003c,16'h000a,16'h001f,16'h0000,-16'h000d,-16'h0010,-16'h000c,-16'h002f,16'h002f,16'h0026,-16'h00b7,16'h0025,16'h003f,-16'h002c,16'h001b,16'h0047,16'h0023,-16'h0028,-16'h003c,16'h001a,16'h000e,16'h002a,16'h000a,-16'h0030,-16'h005d,-16'h000b,16'h0017,16'h001f,-16'h003d,16'h0031,-16'h0047,-16'h002b,-16'h004a,-16'h0016,16'h0024,-16'h0029,16'h0079,16'h007b,-16'h000c,16'h0063,16'h004d,16'h0023,16'h002d,-16'h000e,16'h003c,16'h0043,-16'h0004,-16'h005a,-16'h0031,16'h005e,-16'h0002,16'h000e,-16'h0007,-16'h0009,-16'h000c,16'h0033,16'h0005,16'h004a,16'h0017,16'h004f,16'h0028,-16'h001b,-16'h0002,16'h0030,16'h0009,16'h0024,16'h0015,16'h0007,16'h0005,16'h0031,16'h0002,-16'h000f,16'h0029,16'h0034,-16'h00c2,16'h0032,16'h002e,-16'h0008,16'h003d,16'h005e,16'h000f,16'h0000,-16'h0014,16'h0025,16'h0002,16'h0028,16'h0005,-16'h002b,-16'h004d,16'h0007,16'h0007,-16'h0013,-16'h002d,16'h004c,-16'h0020,-16'h0028,-16'h005c,-16'h0032,16'h001c,-16'h0039,16'h008a,16'h0049,-16'h0002,16'h0048,16'h0089,16'h000f,16'h0058,16'h0000,16'h003a,16'h0033,-16'h0009,-16'h004e,-16'h0014,16'h0066,-16'h001b,16'h0017,16'h0001,-16'h0023,16'h0013,16'h0000,16'h000b,16'h0003,-16'h0017,16'h0059,16'h003f,-16'h000e,16'h000f,16'h0037,16'h0026,16'h0020,16'h0029,16'h002c,-16'h001b,16'h004c,-16'h0019,-16'h0031,16'h000a,16'h0034,-16'h0097,-16'h001e,16'h001d,-16'h0010,16'h002e,16'h006c,16'h001a,16'h0016,-16'h000e,16'h0024,-16'h0005,16'h0025,16'h0012,-16'h002f,-16'h003d,16'h0015,16'h0014,-16'h000d,-16'h002a,16'h0030,-16'h0013,-16'h0034,-16'h0048,-16'h0002,16'h000f,-16'h000e,16'h006e,-16'h000d,16'h0002,16'h0032,16'h0080,16'h000d,16'h005e,-16'h000d,16'h003f,16'h003b,-16'h0019,-16'h001c,16'h0016,16'h0064,-16'h0039,16'h0011,16'h0023,-16'h0017,16'h002f,-16'h0002,16'h001d,-16'h0018,-16'h0022,16'h0061,16'h0035,16'h0006,16'h0012,16'h0008,-16'h000f,-16'h0051,16'h0029,16'h000c,-16'h0014,16'h001d,16'h003e,-16'h0063,16'h0001,16'h0002,16'h0027,16'h001d,-16'h0014,-16'h0083,16'h0029,16'h0063,16'h0008,16'h000e,16'h0013,16'h0023,-16'h0022,-16'h0005,16'h0050,16'h0032,-16'h005a,16'h003a,-16'h000d,16'h0010,16'h000c,16'h0006,-16'h0041,-16'h004b,-16'h0024,-16'h0033,-16'h000f,16'h0008,16'h005a,16'h002f,-16'h000e,16'h0044,-16'h0033,16'h0066,16'h0030,16'h0029,-16'h0029,-16'h0035,16'h003e,16'h0008,16'h0027,-16'h0034,16'h0000,-16'h003b,-16'h0033,16'h0015,16'h004f,-16'h0066,16'h0032,-16'h0019,16'h003c,-16'h000c,-16'h0016,-16'h0038,-16'h0031,-16'h0030,-16'h002a,-16'h0017,16'h003e,16'h002b,-16'h000c,-16'h000d,16'h002c,-16'h009a,16'h0049,-16'h0004,-16'h0009,16'h003a,-16'h0003,-16'h0058,16'h0050,16'h005b,16'h001c,16'h001f,-16'h000d,16'h0011,-16'h001f,-16'h0020,16'h00b4,16'h003f,-16'h0047,16'h0031,16'h0000,16'h0005,16'h0022,16'h0017,-16'h0048,-16'h0014,-16'h0026,16'h000a,16'h0002,16'h002a,16'h0070,16'h0034,-16'h002c,16'h0033,-16'h002d,16'h005f,16'h0023,16'h0034,-16'h0030,-16'h0030,16'h0023,-16'h0004,-16'h0005,-16'h0050,-16'h005e,-16'h0039,-16'h0001,-16'h002f,16'h005c,-16'h002a,16'h001d,-16'h0001,-16'h0011,-16'h0028,-16'h0037,-16'h0042,-16'h0035,-16'h0003,-16'h002b,-16'h000d,16'h006c,-16'h0012,-16'h002e,-16'h0027,16'h003b,-16'h00a1,16'h0036,16'h002d,-16'h002d,16'h003a,16'h000a,-16'h0042,16'h0043,16'h005c,16'h0028,16'h000d,-16'h0010,16'h001f,-16'h0032,-16'h004c,16'h00b5,16'h001e,-16'h003d,16'h003e,-16'h0003,-16'h0009,16'h001d,16'h001b,-16'h003f,-16'h000c,-16'h000c,16'h0017,-16'h0038,16'h0014,16'h008e,16'h0004,-16'h0041,16'h0053,-16'h0025,16'h007c,16'h0033,16'h0028,-16'h0034,-16'h0007,16'h005b,-16'h004e,16'h0029,-16'h006b,-16'h006c,-16'h0050,-16'h001a,-16'h002e,16'h0056,-16'h0021,16'h002a,16'h0012,-16'h0018,-16'h0021,-16'h0019,-16'h0040,-16'h002d,16'h0038,-16'h005f,-16'h0004,16'h006f,-16'h0031,-16'h0034,16'h0004,16'h0040,-16'h0082,16'h001c,16'h0024,-16'h0058,16'h0069,16'h0019,16'h0013,16'h0035,16'h0021,16'h0009,16'h0010,-16'h0023,16'h002f,-16'h0023,-16'h0046,16'h00a3,16'h001b,-16'h0017,16'h003c,16'h0003,-16'h0014,-16'h0014,16'h000f,-16'h0009,-16'h0002,-16'h0034,16'h002e,-16'h0055,16'h0017,16'h0089,16'h000f,-16'h0028,16'h0045,-16'h0029,16'h004f,16'h003d,16'h001f,-16'h0034,16'h0016,16'h002a,-16'h002e,16'h0048,-16'h0091,-16'h00a3,-16'h003b,-16'h001a,-16'h0040,16'h004d,16'h0008,16'h0036,16'h000b,-16'h0024,16'h0001,-16'h0003,-16'h0022,-16'h000d,16'h0041,-16'h00a9,16'h0003,16'h00a6,-16'h0041,-16'h0022,16'h0014,16'h0018,-16'h006a,16'h0029,16'h000f,-16'h009d,16'h0059,16'h0012,16'h000f,16'h0037,-16'h0024,16'h0017,16'h000a,-16'h0016,16'h0032,-16'h000e,-16'h004d,16'h0062,16'h001a,16'h0000,16'h002b,-16'h0027,-16'h0001,16'h0000,16'h0010,-16'h000e,16'h000b,-16'h0053,16'h0018,-16'h0046,16'h0014,16'h0085,-16'h0011,-16'h0015,16'h0048,-16'h0008,16'h0030,16'h0024,16'h0044,-16'h0038,16'h0021,16'h0014,-16'h0042,16'h004d,-16'h00c0,-16'h0083,-16'h0055,-16'h0009,-16'h0023,16'h0047,16'h0020,16'h0033,16'h0017,16'h000c,-16'h0028,-16'h0029,-16'h0016,-16'h001b,16'h003c,-16'h00bd,16'h000c,16'h00a7,-16'h003c,-16'h0004,16'h0010,16'h0017,-16'h002a,16'h000f,-16'h000b,-16'h00b9,16'h005a,16'h0001,16'h0041,16'h0014,-16'h0077,16'h0019,-16'h0002,-16'h0004,16'h0038,16'h0008,-16'h004e,-16'h000f,16'h0011,-16'h0012,16'h002e,-16'h0022,-16'h0007,16'h0000,16'h0018,16'h002f,16'h0012,-16'h0075,16'h002a,-16'h003e,16'h002e,16'h0094,-16'h001f,-16'h0001,16'h002b,16'h0028,16'h0034,16'h0031,16'h004f,-16'h002a,16'h0005,-16'h0007,-16'h005f,16'h005e,-16'h00cb,-16'h001f,-16'h0065,16'h001f,-16'h001d,16'h0070,16'h003c,16'h002c,16'h001d,-16'h000b,16'h000d,-16'h0007,-16'h001d,-16'h000c,16'h005e,-16'h00c8,16'h0042,16'h0096,-16'h0015,-16'h000f,16'h0030,-16'h0011,-16'h001d,-16'h000b,-16'h002c,-16'h00b3,16'h004d,16'h000b,16'h0025,16'h001e,-16'h006a,16'h0007,-16'h0014,-16'h0022,16'h0028,16'h000d,-16'h005a,-16'h0084,16'h0027,-16'h0020,16'h003c,-16'h0021,-16'h0015,-16'h0005,16'h0000,16'h0042,16'h0025,-16'h0067,-16'h0003,16'h0000,-16'h0003,16'h008d,-16'h003f,-16'h000b,16'h0054,16'h002a,-16'h000e,16'h0013,16'h004c,-16'h003a,-16'h000b,-16'h001b,-16'h0089,16'h0030,-16'h00b8,-16'h0006,-16'h005e,16'h0032,16'h0005,16'h0054,16'h0047,16'h0023,16'h0041,-16'h000b,16'h0004,-16'h0002,-16'h0027,16'h0001,16'h0057,-16'h006e,16'h004a,16'h00a6,-16'h000a,-16'h000f,16'h0008,-16'h002d,16'h0000,-16'h000a,-16'h0021,-16'h0098,16'h0030,-16'h001f,16'h0007,-16'h0003,-16'h0042,16'h0011,-16'h000d,-16'h001b,16'h002a,16'h000e,-16'h0079,-16'h0113,16'h0021,-16'h0005,16'h002d,-16'h0008,-16'h000a,16'h0012,16'h0027,16'h003c,16'h0009,-16'h004e,16'h0005,16'h0022,16'h0010,16'h00a2,-16'h003b,-16'h0014,16'h0051,16'h0024,16'h0021,16'h0034,16'h0029,-16'h005b,-16'h0019,16'h0002,-16'h00a0,-16'h0007,-16'h004a,-16'h0024,-16'h0068,16'h004b,16'h000b,16'h0034,16'h0042,16'h0013,16'h003a,16'h0004,16'h0000,16'h0012,-16'h001f,16'h0005,16'h0061,-16'h0042,16'h0044,16'h00a4,-16'h0016,-16'h0013,-16'h0005,-16'h0024,16'h000f,-16'h0015,-16'h0049,-16'h006d,16'h002f,-16'h0012,-16'h000c,-16'h0006,-16'h0067,-16'h0002,16'h0002,-16'h0005,16'h0027,16'h000c,-16'h0061,-16'h0134,16'h0045,16'h000b,16'h001d,-16'h0014,-16'h0010,16'h0005,-16'h0004,16'h0062,-16'h0003,-16'h003d,-16'h000f,16'h0042,-16'h002f,16'h00b7,-16'h0033,-16'h000f,16'h0057,16'h000f,16'h0010,16'h003d,16'h000e,-16'h0067,-16'h000f,-16'h003b,-16'h00a3,-16'h001b,-16'h002b,-16'h0013,-16'h0057,16'h0026,16'h0013,16'h001b,16'h0063,16'h0000,16'h0033,16'h0001,16'h0030,16'h0005,-16'h0039,-16'h001c,16'h001a,-16'h0016,16'h0006,16'h00a5,-16'h0021,-16'h0005,-16'h0028,-16'h003e,16'h0006,-16'h000d,-16'h0033,-16'h005b,16'h0002,16'h000f,-16'h000e,16'h0028,-16'h0066,-16'h000a,-16'h000b,16'h000a,-16'h0008,16'h002f,-16'h006a,-16'h0123,16'h0011,-16'h0009,16'h000b,16'h0000,-16'h0016,16'h000f,-16'h0019,16'h006b,-16'h0001,-16'h0023,16'h0011,16'h0054,-16'h0016,16'h00a0,-16'h001d,-16'h001b,16'h0060,16'h000a,16'h0019,16'h0012,-16'h0003,-16'h009f,-16'h002f,-16'h0032,-16'h0096,-16'h0028,16'h0014,-16'h0016,-16'h0052,16'h001c,16'h0002,16'h000e,16'h0035,16'h0002,16'h001f,-16'h0015,16'h0004,-16'h0006,-16'h0039,-16'h0024,16'h0016,-16'h0008,16'h0000,16'h00aa,-16'h0015,16'h0000,-16'h0015,-16'h000c,16'h002c,16'h0000,-16'h0036,-16'h0036,-16'h001b,-16'h0008,-16'h0017,16'h0015,-16'h0057,-16'h001f,-16'h0015,-16'h0019,16'h0012,16'h0035,-16'h0046,-16'h00e5,16'h0021,16'h0005,16'h001c,16'h000b,-16'h0001,16'h001a,-16'h002a,16'h004a,-16'h0019,-16'h0023,-16'h000a,16'h006f,-16'h0003,16'h0097,16'h0009,-16'h001e,16'h0060,16'h0007,16'h000b,16'h0037,-16'h0015,-16'h00e8,-16'h003d,-16'h0020,-16'h00a7,-16'h0029,16'h001a,-16'h001d,-16'h002d,16'h001a,-16'h000f,16'h0006,-16'h002b,16'h0005,16'h002c,-16'h0024,16'h001e,-16'h0006,-16'h004e,-16'h0002,16'h0003,16'h002c,-16'h0035,16'h0082,-16'h0013,16'h003f,-16'h0018,16'h000d,16'h0057,16'h0011,-16'h0033,-16'h003f,-16'h0019,-16'h0003,-16'h0027,16'h0006,-16'h0043,-16'h0022,-16'h002b,16'h0004,16'h0008,16'h0053,-16'h004b,-16'h009c,16'h0021,-16'h001f,16'h0014,16'h0038,-16'h0011,16'h0008,-16'h003b,16'h004d,-16'h001b,-16'h0020,16'h0003,16'h0052,16'h001e,16'h009e,-16'h0005,-16'h001a,16'h0069,16'h0014,16'h000c,16'h0022,-16'h000d,-16'h0123,-16'h006d,-16'h002b,-16'h009c,-16'h0031,-16'h0023,-16'h0010,-16'h002a,16'h0018,16'h001d,16'h0007,-16'h0056,-16'h0018,16'h0028,-16'h0014,16'h0003,-16'h000d,-16'h002d,-16'h0007,16'h001e,16'h0012,-16'h0038,16'h0077,16'h0009,16'h0037,-16'h0024,16'h000c,16'h0066,16'h001e,16'h000e,-16'h003b,-16'h004c,-16'h0005,16'h0026,-16'h0004,-16'h001e,16'h0003,-16'h000c,-16'h000b,16'h0011,16'h0050,-16'h006d,-16'h003b,16'h000b,16'h0007,-16'h0011,16'h0039,-16'h000a,-16'h0010,-16'h0016,16'h002b,-16'h0014,-16'h0006,16'h0015,16'h002b,-16'h0006,16'h00a0,16'h002a,-16'h000f,16'h004f,16'h0009,-16'h0004,16'h0038,16'h0002,-16'h0134,-16'h00a5,-16'h0012,-16'h00a4,-16'h0042,16'h0017,-16'h001d,-16'h001c,16'h000d,16'h000f,-16'h001a,-16'h0074,-16'h0018,16'h0047,-16'h000b,-16'h000a,16'h0005,-16'h0021,16'h0000,16'h000d,16'h0012,-16'h004f,16'h008c,-16'h0001,16'h003c,-16'h0020,16'h0009,16'h008d,16'h000d,-16'h0006,-16'h0020,-16'h0038,16'h0005,16'h0062,16'h002c,-16'h001b,16'h0005,-16'h0034,-16'h0015,16'h0011,16'h0043,-16'h004f,16'h0016,-16'h000b,16'h0019,16'h0027,16'h002e,-16'h0034,-16'h0019,-16'h0002,16'h0020,-16'h0002,-16'h000c,-16'h0006,-16'h0009,-16'h0022,16'h00bc,16'h0027,-16'h0026,16'h007e,16'h0007,-16'h001c,16'h003a,16'h0013,-16'h00ff,-16'h00a8,-16'h0003,-16'h00a4,-16'h005a,16'h0002,-16'h0002,-16'h0022,16'h0001,16'h0038,-16'h000b,-16'h0051,-16'h001d,16'h0031,16'h0010,-16'h000e,-16'h000b,-16'h002f,16'h0008,16'h000f,16'h0028,-16'h0058,16'h0081,-16'h0006,16'h001c,-16'h000e,16'h0012,16'h0083,16'h000e,16'h0019,16'h0035,-16'h0052,16'h0021,16'h0069,16'h003a,16'h0011,-16'h0002,-16'h0001,-16'h0011,16'h0021,16'h0033,16'h0003,16'h0049,-16'h0011,16'h002b,16'h0020,16'h0002,-16'h000e,-16'h0030,16'h000a,16'h002a,16'h0003,16'h0000,16'h001e,-16'h0031,-16'h000c,16'h00b6,16'h0049,-16'h0022,16'h008b,16'h003c,-16'h0042,16'h005a,-16'h0009,-16'h00e1,-16'h00a1,16'h0020,-16'h00b6,-16'h0088,-16'h0003,-16'h0010,-16'h0016,16'h0001,16'h0029,-16'h000f,-16'h0031,16'h0022,16'h002f,16'h000a,-16'h0025,16'h0017,-16'h0033,-16'h0021,16'h0010,16'h0019,-16'h0031,16'h006c,-16'h001a,-16'h0003,-16'h000b,16'h0002,16'h0081,16'h001c,16'h001a,16'h0085,-16'h003a,-16'h0008,16'h0044,16'h0045,16'h0007,-16'h0005,-16'h0003,-16'h000b,16'h0018,16'h0011,16'h002a,16'h003b,-16'h000a,16'h0020,16'h0006,16'h0011,16'h000a,-16'h0028,16'h0003,16'h0027,16'h000f,-16'h000e,16'h0003,-16'h001e,16'h0018,16'h0090,16'h003e,-16'h0043,16'h009d,16'h0022,-16'h002d,16'h0024,-16'h0018,-16'h00e6,-16'h00c6,16'h0009,-16'h00a3,-16'h005d,16'h0024,16'h0002,16'h0000,16'h000f,16'h0037,16'h0010,-16'h000c,16'h0015,-16'h0004,16'h0006,-16'h0015,16'h0007,-16'h0020,-16'h001d,16'h0000,16'h0028,16'h0003,16'h0078,-16'h001a,-16'h0038,16'h0003,16'h0010,16'h0086,16'h0014,16'h0003,16'h005f,-16'h0021,-16'h000d,-16'h0023,16'h0054,16'h0012,-16'h0009,-16'h001c,16'h000f,16'h001b,-16'h0019,16'h004f,16'h0042,-16'h0017,-16'h0011,16'h0030,16'h0004,16'h0018,-16'h0054,16'h0022,16'h0036,-16'h0010,-16'h0026,16'h0018,16'h0000,16'h002e,16'h0078,16'h0049,-16'h0036,16'h0094,16'h0032,-16'h0044,-16'h0002,-16'h003d,-16'h009d,-16'h00d4,16'h0028,-16'h009a,-16'h0065,16'h0009,16'h0005,-16'h000d,16'h0030,16'h0046,16'h001a,-16'h0019,16'h003e,-16'h001a,16'h000d,-16'h003e,16'h0012,-16'h001a,-16'h0023,16'h0002,16'h0020,16'h000a,16'h0061,-16'h001c,-16'h0056,16'h0008,16'h0014,16'h0053,16'h0014,16'h0009,16'h005b,-16'h0017,-16'h0023,-16'h006a,16'h0040,16'h0036,-16'h0013,16'h0000,16'h000d,16'h001f,-16'h0087,16'h0059,16'h0027,-16'h0033,-16'h005d,16'h0016,-16'h001b,16'h000f,-16'h003f,16'h0010,16'h0044,16'h001a,-16'h0026,16'h001e,-16'h0001,16'h003f,16'h0077,16'h0039,-16'h003b,16'h0097,16'h000d,-16'h003a,-16'h001a,-16'h006f,-16'h0067,-16'h009f,16'h001e,-16'h009b,-16'h0067,-16'h0015,-16'h000a,-16'h0006,16'h000c,16'h0049,16'h0012,16'h0034,16'h0026,-16'h001c,16'h000c,-16'h0031,16'h001f,16'h0000,-16'h0004,16'h0004,16'h0007,16'h0022,16'h006a,-16'h0012,-16'h0045,-16'h000f,-16'h0007,16'h0043,-16'h0024,16'h0006,16'h003a,16'h0026,-16'h0013,-16'h0027,16'h0024,16'h000c,-16'h0032,16'h0023,16'h0015,16'h0020,-16'h013d,16'h005b,16'h000f,-16'h0024,-16'h0048,16'h0009,-16'h003f,-16'h0016,-16'h0013,16'h0029,16'h000a,16'h0008,-16'h0032,16'h002d,-16'h0019,16'h0047,16'h0069,-16'h0006,-16'h001d,16'h0074,16'h0012,-16'h001d,-16'h0027,-16'h00be,-16'h0046,-16'h00b5,16'h003f,-16'h009f,-16'h0066,16'h000e,16'h0010,16'h000d,16'h0002,16'h0053,16'h0016,16'h0066,16'h0040,-16'h003b,16'h0038,-16'h0025,16'h0017,-16'h0003,16'h000c,16'h001c,16'h0025,16'h0047,16'h007e,-16'h0007,-16'h000f,-16'h0037,16'h0012,16'h0004,-16'h001e,-16'h000c,16'h0039,16'h0048,-16'h002a,-16'h000f,-16'h0007,16'h0036,-16'h0059,-16'h0001,16'h0023,16'h001d,-16'h01a1,16'h0067,16'h002a,-16'h0012,-16'h0028,16'h0008,-16'h0006,16'h0007,16'h003a,16'h000d,-16'h0018,16'h000a,-16'h0048,16'h0026,-16'h004d,16'h0040,16'h0065,-16'h007c,-16'h0045,16'h0088,16'h0008,16'h0020,-16'h001a,-16'h00e2,16'h000d,-16'h008e,16'h0013,-16'h00cd,-16'h005f,16'h000f,16'h0018,16'h0007,16'h001f,16'h0046,16'h002b,16'h0066,16'h0035,-16'h002c,16'h003a,-16'h0016,-16'h0007,-16'h0001,16'h004f,16'h0011,16'h0053,16'h0032,16'h0070,-16'h0003,16'h0007,-16'h0024,16'h0007,-16'h0027,-16'h000e,-16'h000c,16'h0025,16'h006e,-16'h0023,16'h0007,-16'h005b,16'h002e,-16'h0054,16'h0017,16'h001f,16'h0016,-16'h0141,16'h0068,16'h001d,16'h0004,16'h000b,16'h001b,16'h000a,-16'h001c,16'h0055,-16'h000d,-16'h0081,-16'h000e,-16'h0032,16'h001b,-16'h0055,16'h001b,16'h002a,-16'h0041,-16'h0027,16'h0099,16'h0003,16'h0025,-16'h003b,-16'h0115,16'h0053,-16'h00a3,16'h001a,-16'h00a1,-16'h0078,16'h001e,16'h000b,16'h000c,16'h000c,16'h0026,16'h003d,16'h0054,16'h004d,-16'h0031,16'h0050,16'h0010,-16'h0004,16'h0003,16'h0041,16'h000a,16'h0064,16'h0024,16'h0052,16'h0017,-16'h002d,-16'h0019,-16'h0019,-16'h007a,16'h0023,-16'h0007,16'h000d,16'h0062,-16'h0003,-16'h0017,-16'h0125,16'h0031,-16'h0041,16'h000e,16'h001b,16'h001c,-16'h0095,16'h0036,16'h002e,16'h0035,-16'h000e,16'h0019,16'h001c,-16'h000a,16'h002f,-16'h0005,-16'h00a9,-16'h0009,-16'h0053,16'h0014,-16'h0038,-16'h0033,16'h0016,16'h000d,-16'h001d,16'h008c,16'h0008,16'h004a,-16'h0037,-16'h00fa,16'h0061,-16'h008b,16'h000a,-16'h0083,-16'h006a,16'h0015,16'h000c,16'h0014,16'h0015,16'h001f,16'h0015,16'h0034,16'h005f,-16'h0008,16'h003c,16'h0031,16'h001d,-16'h0004,16'h0074,16'h000a,16'h006a,16'h0020,16'h0038,16'h000b,16'h0000,16'h0013,16'h0012,-16'h0089,16'h0025,-16'h0009,-16'h0020,16'h006e,16'h002b,-16'h0014,-16'h014c,16'h004d,-16'h0003,16'h0010,16'h0007,16'h0061,-16'h0060,16'h003c,16'h0029,16'h0020,16'h0011,16'h0015,16'h0034,-16'h0003,16'h0015,-16'h002c,-16'h0095,-16'h0010,-16'h0042,-16'h0012,-16'h001e,-16'h0053,16'h0043,16'h0052,-16'h0020,16'h00ac,16'h0017,16'h002d,-16'h0025,-16'h00cb,16'h0070,-16'h0049,-16'h0049,-16'h006b,-16'h0020,16'h002a,-16'h000f,16'h001f,16'h002a,-16'h0009,16'h000f,16'h0012,16'h006f,16'h0011,16'h0067,16'h005a,16'h0006,-16'h0029,16'h0055,-16'h0001,16'h0062,16'h001f,16'h0041,16'h001e,-16'h0002,16'h000d,16'h0015,-16'h0066,16'h001b,16'h0023,-16'h0084,16'h0046,16'h0045,-16'h0020,-16'h00e8,16'h0048,16'h0019,16'h000e,-16'h000f,16'h0030,-16'h004d,16'h0030,16'h0036,-16'h0004,-16'h0038,-16'h001c,16'h004e,-16'h000b,-16'h001e,-16'h001a,-16'h00a4,-16'h000d,-16'h0040,16'h000d,-16'h0001,-16'h0041,16'h002f,16'h00a2,-16'h003b,16'h009d,16'h0054,16'h002c,-16'h001f,-16'h0081,16'h0084,-16'h0006,-16'h0047,-16'h0081,16'h0002,16'h0042,-16'h0023,16'h0026,16'h0020,-16'h0019,16'h0019,-16'h000d,16'h0059,16'h004c,16'h005d,16'h0054,-16'h0005,-16'h0036,16'h003f,16'h000b,16'h005d,16'h0020,16'h001a,16'h0048,-16'h002b,16'h001c,-16'h000d,-16'h0063,16'h0028,16'h001d,-16'h00b8,16'h0029,16'h002d,-16'h0017,-16'h004d,16'h005f,16'h003f,-16'h0007,-16'h0020,16'h0011,-16'h000d,16'h0012,16'h0004,-16'h0039,-16'h0018,-16'h0017,16'h0037,-16'h0007,-16'h002f,-16'h0034,-16'h0054,-16'h0008,-16'h0059,-16'h0012,16'h0017,-16'h002f,16'h004b,16'h009b,-16'h0026,16'h0094,16'h003b,16'h0026,-16'h0021,-16'h0046,16'h006e,16'h003f,-16'h003a,-16'h007f,-16'h000e,16'h005d,-16'h000f,16'h000e,16'h0018,-16'h0062,16'h0036,-16'h0002,16'h0039,16'h0057,16'h0058,16'h007f,-16'h0001,-16'h0020,16'h0028,16'h0025,16'h0056,16'h0037,16'h0017,16'h0032,-16'h0002,16'h0016,-16'h000f,-16'h005f,16'h0026,16'h0036,-16'h00fc,16'h0034,16'h0021,-16'h001f,16'h0030,16'h005d,16'h0035,16'h0007,-16'h002f,16'h0027,-16'h0019,16'h000c,16'h000c,-16'h0052,-16'h0044,16'h0008,16'h0027,16'h000f,-16'h003f,16'h002d,-16'h0030,-16'h0026,-16'h0064,-16'h000e,-16'h000c,-16'h0022,16'h0066,16'h0079,-16'h0017,16'h0090,16'h0043,16'h001e,16'h000d,-16'h0032,16'h005a,16'h0055,-16'h0025,-16'h0072,16'h0003,16'h0053,-16'h0019,-16'h0010,-16'h000d,-16'h0043,16'h0037,16'h001f,16'h000c,16'h0037,16'h0009,16'h005f,16'h0030,-16'h0025,16'h0026,16'h0040,16'h0033,16'h0025,16'h0022,16'h0029,-16'h0007,16'h0029,16'h0007,-16'h003c,16'h002f,16'h0041,-16'h00e1,16'h003c,16'h0042,-16'h0024,16'h0033,16'h0042,16'h004b,-16'h0023,-16'h0019,16'h000f,-16'h000a,16'h0000,-16'h0001,-16'h0059,-16'h0047,16'h0005,16'h0009,-16'h001e,-16'h003f,16'h0043,-16'h002b,-16'h0020,-16'h0072,-16'h000a,-16'h000f,-16'h0019,16'h009e,16'h003c,16'h0009,16'h0066,16'h0051,16'h0032,16'h0033,-16'h0010,16'h005f,16'h0041,16'h0003,-16'h0065,16'h0002,16'h0055,-16'h000c,-16'h000f,-16'h0002,-16'h0036,16'h0019,16'h0004,16'h000c,16'h0036,-16'h001d,16'h0059,16'h0029,-16'h0019,16'h0015,16'h002a,16'h0035,16'h0031,16'h0031,16'h001b,-16'h000d,16'h002c,-16'h000c,-16'h0049,16'h001a,16'h0019,-16'h00ba,16'h0009,16'h0032,16'h000c,16'h0040,16'h004e,16'h0037,16'h0011,16'h0006,16'h0030,16'h0010,-16'h0001,-16'h001a,-16'h003f,-16'h004c,16'h0033,16'h0012,16'h0007,-16'h0033,16'h0028,-16'h001b,-16'h001a,-16'h0055,-16'h000a,16'h000a,-16'h0019,16'h0093,16'h001b,16'h0006,16'h002b,16'h006f,16'h0015,16'h0042,-16'h001c,16'h005e,16'h0046,16'h000d,-16'h0050,16'h0031,16'h0070,-16'h0043,16'h0004,16'h001e,-16'h0022,16'h001c,-16'h0003,16'h000f,16'h0006,-16'h004e,16'h0070,16'h0040,-16'h0005,16'h0005,-16'h000f,-16'h002d,-16'h0034,16'h003d,16'h0005,-16'h0020,16'h000e,16'h008d,-16'h006e,16'h0030,16'h0020,16'h0013,16'h0011,-16'h0026,-16'h007a,16'h0041,16'h0089,-16'h0002,16'h0003,-16'h0001,16'h002f,-16'h0022,-16'h0003,16'h0072,16'h0038,-16'h002b,16'h005a,16'h0010,16'h0005,16'h0007,-16'h0008,-16'h0060,-16'h003e,-16'h001d,-16'h0004,-16'h0011,16'h0018,16'h004c,16'h002b,16'h0001,16'h0040,-16'h002e,16'h0079,16'h0005,16'h0042,-16'h0013,-16'h0041,16'h003b,-16'h0029,16'h002a,-16'h005a,-16'h001d,-16'h0045,-16'h002b,16'h0002,16'h005e,-16'h0040,16'h002b,-16'h0035,16'h0020,-16'h0023,-16'h000a,-16'h0041,-16'h0029,16'h0000,-16'h003e,-16'h002c,16'h004f,-16'h0016,-16'h0018,16'h0012,16'h0085,-16'h00ba,16'h0060,16'h001a,16'h0003,16'h0037,-16'h000c,-16'h0060,16'h0037,16'h0059,16'h001c,16'h0011,-16'h000d,16'h0032,-16'h003a,-16'h003c,16'h00b4,16'h0025,-16'h002c,16'h0036,16'h0009,-16'h0002,16'h001b,16'h0010,-16'h003b,-16'h0034,-16'h0004,16'h0008,-16'h0015,16'h000d,16'h0084,16'h005b,16'h0010,16'h002d,-16'h0023,16'h0073,16'h0053,16'h003b,-16'h0029,-16'h0007,16'h001a,-16'h000d,16'h003c,-16'h0072,-16'h0061,-16'h002d,-16'h0027,-16'h0021,16'h0053,-16'h0026,16'h0057,-16'h001a,16'h0001,-16'h0010,-16'h0005,-16'h005c,-16'h0032,16'h000d,-16'h006e,-16'h001d,16'h0063,-16'h0017,-16'h0031,-16'h000d,16'h0040,-16'h00b1,16'h0041,16'h002f,-16'h0030,16'h0063,-16'h0005,-16'h004b,16'h0030,16'h0036,16'h0045,16'h000a,-16'h002f,16'h0047,-16'h004c,-16'h003c,16'h00c3,16'h002c,-16'h000c,16'h0032,-16'h0001,-16'h001b,16'h000b,16'h0018,-16'h002e,-16'h000f,-16'h0009,16'h0009,-16'h0044,16'h001e,16'h0071,16'h0019,-16'h0012,16'h002e,-16'h005f,16'h0064,16'h0036,16'h001d,-16'h0032,-16'h0005,16'h0042,-16'h0021,16'h002a,-16'h00ba,-16'h0089,-16'h0046,-16'h001a,-16'h0020,16'h004a,-16'h002c,16'h0052,-16'h0004,16'h0007,16'h0000,16'h0000,-16'h003f,-16'h0008,16'h003c,-16'h009d,-16'h0034,16'h009f,-16'h0033,-16'h0042,16'h001e,16'h003b,-16'h0086,16'h0014,16'h0053,-16'h008a,16'h0050,16'h000f,16'h0012,16'h0031,16'h0004,16'h0021,16'h0008,-16'h0037,16'h0041,-16'h0030,-16'h004e,16'h0066,16'h0025,-16'h0028,16'h0052,-16'h001c,16'h0007,-16'h0024,16'h000c,16'h0002,-16'h001e,-16'h0024,16'h0015,-16'h004b,-16'h0011,16'h0086,-16'h0003,16'h0028,16'h0038,-16'h0048,16'h002b,16'h0023,16'h002a,-16'h0038,16'h0004,16'h001b,-16'h0018,16'h005c,-16'h00c7,-16'h00a7,-16'h004d,16'h0008,-16'h0032,16'h006e,16'h0004,16'h0057,16'h0034,16'h0018,16'h0008,-16'h0029,-16'h0034,-16'h0038,16'h005e,-16'h00d6,-16'h0015,16'h00a6,-16'h004d,-16'h0025,16'h0034,16'h0017,-16'h0069,16'h0013,16'h0015,-16'h00d2,16'h0081,16'h001c,16'h0049,16'h0035,-16'h0025,16'h002d,-16'h0002,-16'h002a,16'h002b,-16'h0006,-16'h0042,16'h001b,16'h0018,-16'h001e,16'h0052,-16'h0023,16'h001d,-16'h0011,16'h0006,16'h0012,16'h0004,-16'h0047,16'h001e,-16'h004f,16'h0018,16'h00ab,16'h000a,16'h005d,16'h0042,16'h0001,16'h001f,16'h0019,16'h0035,-16'h003d,16'h0016,16'h0016,-16'h0054,16'h007f,-16'h00aa,-16'h0077,-16'h004c,16'h001f,-16'h0013,16'h006a,16'h000c,16'h005b,16'h003d,16'h000c,16'h0000,16'h0004,-16'h001b,-16'h0022,16'h006e,-16'h00d1,16'h002a,16'h0083,-16'h003a,-16'h0015,16'h003e,16'h0016,-16'h0013,16'h0004,-16'h0028,-16'h00bb,16'h0075,16'h000e,16'h002b,16'h000c,-16'h0061,16'h0040,-16'h0016,-16'h002f,16'h004d,16'h001d,-16'h0049,-16'h0061,16'h0000,-16'h0023,16'h0059,-16'h003c,16'h0004,-16'h0011,-16'h0007,16'h0051,-16'h0007,-16'h0037,-16'h0010,-16'h002f,16'h0020,16'h00be,-16'h000f,16'h005d,16'h0049,16'h0018,16'h0028,16'h000d,16'h0032,-16'h004d,-16'h0029,16'h001c,-16'h0088,16'h0077,-16'h0092,-16'h000f,-16'h003f,16'h0030,-16'h001e,16'h007c,16'h005a,16'h0046,16'h0050,-16'h0007,16'h0004,16'h0009,-16'h0014,-16'h000c,16'h0071,-16'h0077,16'h0042,16'h0097,-16'h0020,-16'h0025,16'h0025,-16'h0018,-16'h000b,-16'h0012,-16'h0037,-16'h00ce,16'h007b,16'h0010,16'h0005,16'h0005,-16'h0052,16'h0050,-16'h001b,-16'h000f,16'h0038,16'h0001,-16'h0065,-16'h00ed,16'h0026,16'h000f,16'h0049,-16'h0012,-16'h0009,16'h0003,16'h000f,16'h0043,-16'h0035,-16'h0058,16'h0000,16'h0022,16'h001d,16'h00aa,-16'h000e,16'h0053,16'h004d,16'h003f,16'h0026,16'h003e,16'h0014,-16'h0069,-16'h0010,16'h0015,-16'h00a8,16'h0048,-16'h0055,-16'h001d,-16'h0053,16'h0050,-16'h0010,16'h0048,16'h0048,16'h0048,16'h004c,16'h000a,-16'h0019,16'h000f,-16'h000d,-16'h000f,16'h006a,-16'h001d,16'h0039,16'h00a4,-16'h001b,-16'h001b,16'h0017,-16'h000a,16'h0011,-16'h001a,-16'h0028,-16'h007f,16'h0044,-16'h000c,-16'h0021,-16'h0009,-16'h002d,16'h0034,-16'h0019,-16'h0013,16'h0006,16'h0003,-16'h005d,-16'h0131,16'h0044,16'h0000,16'h0047,-16'h0025,-16'h0005,-16'h002f,16'h0002,16'h0066,-16'h0015,-16'h0045,-16'h001b,16'h005a,-16'h0006,16'h009a,-16'h0029,16'h005c,16'h0052,16'h002a,16'h004e,16'h004d,16'h0006,-16'h0050,16'h000b,-16'h0022,-16'h00ae,16'h001d,16'h000c,16'h0003,-16'h004d,16'h002b,-16'h0017,16'h0021,16'h005a,16'h004f,16'h004e,-16'h0013,-16'h000e,-16'h0002,-16'h001e,-16'h0023,16'h0071,16'h0000,16'h0026,16'h00a2,-16'h001f,-16'h0031,16'h0010,-16'h002d,16'h0011,-16'h001c,-16'h001a,-16'h008f,16'h0041,-16'h000f,-16'h0043,16'h001a,-16'h005b,16'h0045,-16'h0002,16'h0010,16'h0030,16'h000b,-16'h008c,-16'h013a,16'h0030,16'h0009,16'h001b,-16'h0025,-16'h001a,-16'h0018,-16'h0010,16'h0061,16'h0000,-16'h000f,-16'h0007,16'h0038,-16'h0030,16'h00b0,-16'h0043,16'h0060,16'h0037,16'h0023,16'h0024,16'h002c,16'h0010,-16'h009a,16'h0010,-16'h001c,-16'h00a4,-16'h0042,16'h0017,-16'h0009,-16'h006e,16'h001f,-16'h000e,-16'h0002,16'h0056,16'h0046,16'h0038,-16'h001f,16'h0000,16'h0020,-16'h0025,-16'h002f,16'h003e,16'h0021,16'h000d,16'h0098,-16'h0027,16'h0000,-16'h000b,-16'h0018,16'h0049,-16'h0009,-16'h003c,-16'h0068,16'h0004,-16'h0006,-16'h003f,16'h0003,-16'h005f,16'h001f,-16'h0012,-16'h0001,16'h0011,16'h0027,-16'h0079,-16'h00cf,16'h0004,-16'h0013,16'h0010,-16'h0022,16'h0003,-16'h0021,-16'h001a,16'h0059,-16'h002a,-16'h0024,16'h000b,16'h006f,-16'h0003,16'h00c3,-16'h0014,16'h0041,16'h004b,16'h001e,16'h002e,16'h0046,-16'h0014,-16'h00f1,16'h0011,-16'h0011,-16'h00bb,-16'h0041,16'h002c,-16'h0016,-16'h0078,16'h000f,-16'h001a,16'h000c,-16'h0002,16'h0012,16'h0050,-16'h001e,-16'h0018,-16'h0009,-16'h001f,-16'h002b,16'h0003,16'h004d,-16'h0027,16'h0073,-16'h0023,16'h0021,-16'h001a,16'h000b,16'h006d,16'h001c,-16'h0038,-16'h004d,-16'h002e,-16'h0019,-16'h000b,16'h0014,-16'h0042,16'h0000,-16'h0021,16'h000b,16'h0018,16'h0044,-16'h006b,-16'h0056,16'h0016,16'h000b,16'h0014,16'h0013,-16'h0020,-16'h0010,-16'h0015,16'h006b,-16'h0019,16'h0013,16'h0021,16'h007d,16'h0015,16'h0096,-16'h0008,16'h0035,16'h0042,16'h0005,16'h002f,16'h0053,16'h0001,-16'h0167,16'h000c,16'h0000,-16'h00e6,-16'h0010,16'h0011,16'h0000,-16'h0070,16'h0015,-16'h0019,16'h0007,-16'h0042,16'h001a,16'h0037,-16'h0025,-16'h001e,16'h000c,-16'h0012,16'h0003,-16'h0005,16'h0034,-16'h003b,16'h005d,16'h0001,16'h0021,-16'h001b,-16'h0003,16'h0070,16'h001a,-16'h002d,-16'h003b,-16'h0024,-16'h0011,16'h001d,-16'h0014,-16'h0037,-16'h000c,-16'h0004,16'h0004,16'h001f,16'h005c,-16'h004f,-16'h0004,16'h0030,-16'h0006,16'h0017,16'h0002,-16'h0012,16'h0022,-16'h0025,16'h0031,16'h0000,-16'h000a,16'h002b,16'h0029,16'h0018,16'h0098,-16'h0015,16'h003f,16'h004b,16'h0012,16'h001e,16'h0031,-16'h0001,-16'h014c,-16'h0012,-16'h0006,-16'h00c8,-16'h0027,-16'h0013,-16'h0013,-16'h0053,16'h0000,16'h0019,16'h0011,-16'h005c,16'h0024,16'h0020,16'h0002,-16'h0026,-16'h0004,-16'h001b,16'h0017,-16'h0026,16'h003f,-16'h0028,16'h0079,16'h000c,16'h002f,-16'h0011,16'h000c,16'h007a,-16'h0005,-16'h0002,-16'h003e,-16'h0057,-16'h000e,16'h005a,16'h0017,-16'h0037,-16'h0004,-16'h0013,-16'h000d,16'h0036,16'h005a,-16'h004a,16'h0040,-16'h0002,-16'h000c,16'h0012,16'h0017,-16'h0006,16'h0020,-16'h001b,16'h0040,-16'h000d,-16'h0019,16'h0010,-16'h000f,-16'h0012,16'h00a0,16'h0006,16'h002c,16'h0064,16'h0026,-16'h0015,16'h0066,16'h0001,-16'h00d9,-16'h001a,16'h0014,-16'h00d5,-16'h0035,-16'h0001,-16'h0008,-16'h0052,-16'h0015,16'h002e,16'h0000,-16'h005d,16'h000a,16'h0025,16'h0005,-16'h0026,-16'h0012,-16'h0029,16'h000f,-16'h0030,16'h0025,-16'h001c,16'h0089,16'h000d,16'h0032,-16'h001c,16'h0000,16'h0088,-16'h0009,-16'h001c,-16'h0019,-16'h0041,16'h000c,16'h0063,16'h0033,-16'h001b,-16'h0001,-16'h002a,-16'h0005,16'h002e,16'h0048,-16'h0002,16'h005c,-16'h0001,16'h0006,16'h0019,16'h000c,-16'h001e,16'h0009,-16'h0015,16'h002f,-16'h0010,-16'h0034,-16'h0004,-16'h001d,-16'h0029,16'h00ad,16'h0023,16'h002c,16'h009e,16'h001f,16'h0003,16'h003a,-16'h000a,-16'h0088,-16'h0042,16'h0019,-16'h00d8,-16'h0058,-16'h000a,-16'h001a,-16'h0067,-16'h0020,16'h003b,16'h000c,-16'h002d,16'h0032,16'h000c,16'h0014,-16'h0023,16'h0004,-16'h000a,16'h0029,16'h0000,16'h0011,-16'h001a,16'h0084,16'h000f,16'h0015,16'h0000,16'h000d,16'h0092,16'h000e,16'h000c,16'h001c,-16'h0037,16'h0004,16'h0052,16'h0049,-16'h0007,16'h001c,-16'h000a,-16'h000c,16'h0025,16'h0053,16'h002e,16'h0054,16'h0019,16'h000d,16'h000e,-16'h0005,-16'h0008,16'h000e,-16'h0009,16'h002d,-16'h0024,-16'h001b,-16'h0018,-16'h0054,-16'h0025,16'h00a6,16'h0024,16'h003a,16'h00a9,16'h002c,-16'h003c,16'h004f,-16'h0016,-16'h0094,-16'h0035,16'h0022,-16'h00c8,-16'h0081,16'h0011,-16'h0013,-16'h007c,16'h000d,16'h0023,-16'h001a,-16'h001e,16'h002a,-16'h000a,-16'h0012,-16'h002e,16'h000b,-16'h0031,-16'h0011,16'h0000,16'h0036,16'h000c,16'h009a,-16'h0013,-16'h000f,-16'h0012,16'h000a,16'h0085,16'h001c,16'h0017,16'h0068,-16'h0034,16'h000c,-16'h0013,16'h003f,16'h0006,16'h003b,-16'h001e,-16'h001c,16'h0034,16'h0028,16'h004c,16'h0072,-16'h000d,16'h0000,16'h0000,16'h000b,16'h0012,-16'h0030,-16'h000e,16'h0023,-16'h0012,-16'h001f,16'h0023,-16'h0021,-16'h000a,16'h008a,16'h0031,16'h0034,16'h00a7,16'h000f,-16'h002d,16'h003b,16'h0024,-16'h0090,-16'h0079,16'h0048,-16'h00c6,-16'h005e,16'h0030,-16'h0023,-16'h004f,16'h000d,16'h0041,-16'h0004,16'h002c,16'h0028,-16'h0001,-16'h0003,-16'h003d,16'h0014,-16'h001f,-16'h0033,16'h000f,16'h002d,16'h0010,16'h0087,-16'h0022,16'h0001,-16'h000e,16'h0015,16'h0060,16'h000b,16'h0005,16'h0063,-16'h0022,-16'h0006,-16'h008a,16'h0070,16'h002d,16'h0022,-16'h0009,16'h000d,16'h0026,-16'h0025,16'h0065,16'h0052,16'h0016,-16'h0023,16'h001e,16'h0006,16'h0009,-16'h003d,-16'h0007,16'h002c,16'h0012,-16'h0021,16'h0010,-16'h0015,16'h0021,16'h008f,16'h004d,16'h0028,16'h00b4,16'h0003,-16'h003e,16'h0012,-16'h000c,-16'h0061,-16'h007e,16'h0042,-16'h00dd,-16'h0061,16'h0021,-16'h001c,-16'h005b,16'h000d,16'h0059,16'h000c,16'h0034,16'h003b,-16'h0026,16'h0004,-16'h003a,16'h0012,-16'h0001,-16'h0016,-16'h0003,16'h0049,16'h001f,16'h0052,-16'h0029,-16'h001e,-16'h000a,16'h0000,16'h0016,-16'h0003,16'h0019,16'h0061,-16'h002a,-16'h0014,-16'h0077,16'h0045,16'h0045,-16'h0010,16'h000e,-16'h0005,16'h002a,-16'h0084,16'h0067,16'h0022,-16'h0014,-16'h004b,16'h0009,-16'h000f,16'h0007,-16'h0054,-16'h0001,16'h0010,16'h002e,-16'h000e,16'h0030,16'h0004,16'h0039,16'h008e,16'h0044,16'h0016,16'h0097,16'h0019,-16'h0048,-16'h0025,-16'h0060,-16'h0031,-16'h0097,16'h0033,-16'h00d6,-16'h0046,16'h0007,-16'h0005,-16'h0040,16'h0032,16'h0063,16'h0010,16'h0047,16'h004c,-16'h0047,16'h0026,-16'h0035,16'h0003,-16'h0018,16'h0002,-16'h0002,16'h0046,16'h0049,16'h0056,-16'h0026,-16'h0016,-16'h0044,16'h0014,-16'h000b,-16'h0015,16'h000c,16'h0069,16'h0027,-16'h0011,-16'h004d,16'h0054,16'h0070,-16'h0010,16'h0012,16'h0013,16'h004a,-16'h0162,16'h0075,16'h000c,-16'h0003,-16'h0043,-16'h001f,-16'h000a,-16'h0027,-16'h001d,-16'h000d,-16'h0013,16'h002f,16'h0001,16'h002e,-16'h0023,16'h0058,16'h0084,-16'h0010,16'h0020,16'h0068,-16'h0018,-16'h0022,-16'h001a,-16'h009f,16'h000b,-16'h009d,16'h004b,-16'h00b2,-16'h0053,16'h0011,-16'h001e,-16'h003b,16'h0018,16'h0068,16'h0014,16'h0051,16'h0042,-16'h0036,16'h0033,-16'h0012,16'h0002,16'h0013,16'h002d,16'h0015,16'h0042,16'h0048,16'h0071,-16'h0032,-16'h0003,-16'h005e,-16'h0019,-16'h002d,-16'h0022,16'h0019,16'h0070,16'h003c,-16'h000f,-16'h002a,16'h0009,16'h0070,-16'h0055,16'h0008,-16'h0002,16'h0048,-16'h01fb,16'h0051,16'h0010,-16'h0004,-16'h002c,16'h0010,16'h000a,-16'h0022,16'h0005,16'h0000,-16'h0042,16'h0000,16'h0012,16'h003c,-16'h0052,16'h0045,16'h006e,-16'h0098,16'h0009,16'h0083,16'h0000,-16'h0009,-16'h002d,-16'h0104,16'h0051,-16'h0090,16'h0039,-16'h00c6,-16'h007a,16'h0016,-16'h000f,-16'h0026,16'h001e,16'h005b,16'h003f,16'h003c,16'h0034,-16'h000a,16'h0037,-16'h000b,16'h0004,16'h0000,16'h005c,-16'h0016,16'h007a,16'h004f,16'h0038,-16'h0006,16'h0013,-16'h0038,-16'h0004,-16'h0064,16'h000b,16'h0019,16'h0042,16'h0054,16'h0024,16'h000e,-16'h0049,16'h0067,-16'h0074,16'h0009,16'h0027,16'h0021,-16'h0159,16'h004c,16'h000e,-16'h001d,-16'h0014,-16'h0001,16'h001f,-16'h001d,16'h006f,16'h0009,-16'h0077,-16'h000e,16'h0010,16'h002c,-16'h0048,16'h0034,16'h0033,-16'h007d,16'h001d,16'h0082,16'h0013,16'h0043,-16'h0031,-16'h0130,16'h0080,-16'h00bd,16'h002e,-16'h00c3,-16'h0067,16'h000e,16'h0012,-16'h0001,16'h0021,16'h005a,16'h003a,16'h0032,16'h004f,16'h000c,16'h0062,16'h0009,16'h0009,16'h0008,16'h0055,-16'h0029,16'h007b,16'h0065,16'h0041,-16'h0010,16'h0029,-16'h004d,16'h0005,-16'h00b0,-16'h000e,16'h0011,16'h0036,16'h0053,16'h0044,16'h0001,-16'h00d4,16'h007b,-16'h0045,16'h0012,16'h0021,16'h0031,-16'h00a2,16'h0016,-16'h0006,16'h0043,-16'h0009,16'h0024,16'h0027,-16'h0017,16'h0060,16'h0002,-16'h00a9,-16'h0017,-16'h000d,16'h0028,-16'h003a,16'h0000,16'h0026,16'h0013,16'h001e,16'h0071,16'h0000,16'h0067,-16'h001f,-16'h0109,16'h007a,-16'h00bc,16'h0016,-16'h00d5,-16'h000d,16'h0002,16'h0019,-16'h0008,16'h000e,16'h0049,16'h003d,16'h0010,16'h0059,16'h000a,16'h0057,16'h0027,16'h001b,-16'h0005,16'h0057,16'h000a,16'h0089,16'h003b,16'h003e,16'h0017,16'h0016,-16'h000e,16'h0001,-16'h00c0,16'h001e,16'h0024,16'h000a,16'h0053,16'h003b,-16'h001c,-16'h0121,16'h0054,-16'h0031,16'h0007,16'h001c,16'h0036,-16'h0078,16'h0010,16'h0022,16'h001c,-16'h000f,-16'h000a,16'h004f,-16'h0027,16'h0023,-16'h0008,-16'h00c0,16'h0001,-16'h003c,16'h0019,-16'h0011,-16'h0042,16'h0033,16'h0085,16'h001a,16'h0081,16'h0023,16'h004a,-16'h0021,-16'h00e9,16'h0096,-16'h0076,-16'h000b,-16'h00a7,16'h000c,16'h0003,16'h0000,-16'h0020,16'h0038,16'h0031,16'h000f,-16'h0019,16'h0087,16'h0013,16'h0060,16'h0057,16'h0025,-16'h0010,16'h0072,16'h0006,16'h0072,16'h0027,16'h0027,16'h002b,16'h002e,16'h0019,16'h001f,-16'h00e0,16'h000a,16'h002d,-16'h003c,16'h005b,16'h001a,16'h0006,-16'h00ce,16'h0075,16'h000b,16'h001b,16'h000b,16'h0053,-16'h002e,16'h0021,16'h0002,-16'h0004,16'h0004,-16'h0022,16'h0034,-16'h003a,-16'h002a,-16'h000f,-16'h0095,-16'h001a,-16'h008a,16'h0020,-16'h0001,-16'h006e,16'h0037,16'h00b8,16'h0004,16'h0077,16'h0025,16'h0030,-16'h0017,-16'h009a,16'h007e,-16'h0047,-16'h0019,-16'h007e,16'h0026,16'h0033,-16'h0024,16'h0007,16'h001b,-16'h0012,16'h000e,-16'h0033,16'h0097,16'h0038,16'h005b,16'h008e,-16'h0016,-16'h0011,16'h0042,16'h0017,16'h0046,16'h002f,16'h0032,16'h0023,16'h003d,16'h0012,-16'h0017,-16'h009d,16'h0014,16'h005e,-16'h009d,16'h0046,16'h0031,-16'h0004,-16'h005d,16'h0066,16'h002e,16'h001b,16'h0015,16'h001f,-16'h001a,16'h002e,-16'h0013,-16'h0013,-16'h0020,-16'h0033,16'h0043,-16'h0023,-16'h0036,-16'h002d,-16'h0070,-16'h0014,-16'h0092,16'h0024,-16'h000f,-16'h004d,16'h0052,16'h00bb,16'h000c,16'h0074,16'h0043,16'h0048,-16'h0022,-16'h005a,16'h0090,-16'h0007,-16'h0042,-16'h0077,16'h0035,16'h003f,-16'h003f,16'h001c,16'h000b,-16'h007a,16'h0025,-16'h0036,16'h0062,16'h002b,16'h0054,16'h0081,-16'h0014,-16'h0024,16'h0032,16'h0017,16'h0047,16'h0034,16'h000a,16'h0039,16'h002e,16'h002e,16'h0012,-16'h0086,16'h001b,16'h005b,-16'h00e1,16'h003e,16'h0033,-16'h000d,16'h001f,16'h0048,16'h0036,16'h0015,-16'h0010,16'h0025,16'h0000,-16'h0003,-16'h0037,-16'h003e,-16'h004a,16'h000d,16'h0025,-16'h0039,-16'h004f,-16'h0012,-16'h0049,-16'h0021,-16'h00b1,16'h0002,-16'h001d,-16'h004c,16'h0079,16'h00a1,16'h0011,16'h0062,16'h0042,16'h0039,16'h0003,-16'h0022,16'h005a,16'h000e,-16'h001c,-16'h0056,16'h0034,16'h0032,16'h0001,16'h0012,-16'h002e,-16'h006a,16'h001c,-16'h0011,16'h003f,16'h004e,16'h003f,16'h0081,16'h0001,-16'h0029,16'h0016,16'h001d,16'h000c,16'h0040,-16'h000b,16'h003b,16'h0011,16'h001a,-16'h000b,-16'h0061,16'h0036,16'h0031,-16'h0115,16'h005f,16'h0038,-16'h0005,16'h0052,16'h0046,16'h005d,-16'h0018,-16'h0031,16'h000c,-16'h0016,-16'h001b,-16'h0033,-16'h004b,-16'h003f,16'h001b,16'h0007,-16'h001e,-16'h0073,16'h003a,-16'h002b,16'h000d,-16'h0090,16'h000c,-16'h0004,-16'h0022,16'h0086,16'h004c,16'h002b,16'h0057,16'h0051,16'h004e,16'h0025,-16'h0018,16'h0046,16'h004e,16'h0009,-16'h0051,16'h001f,16'h003f,-16'h0015,16'h000e,-16'h003e,-16'h0084,16'h0027,16'h000f,16'h000c,16'h0039,-16'h0016,16'h0067,-16'h0004,-16'h0005,-16'h0015,16'h003c,16'h0012,16'h002d,16'h002c,16'h002b,16'h0000,16'h0029,-16'h0002,-16'h0044,16'h003b,16'h0025,-16'h00f3,16'h0027,16'h0045,16'h0014,16'h0054,16'h005b,16'h0054,16'h0010,-16'h0022,16'h001c,-16'h0016,-16'h0014,-16'h0020,-16'h003b,-16'h001d,16'h0013,16'h002a,-16'h0021,-16'h0056,16'h0066,-16'h002f,16'h0008,-16'h0077,16'h0009,16'h0003,16'h0000,16'h0097,16'h0020,16'h000d,16'h0029,16'h0069,16'h002c,16'h0060,-16'h0015,16'h0024,16'h003c,16'h0009,-16'h002b,16'h0047,16'h0071,-16'h0021,16'h0000,-16'h001d,-16'h006d,16'h0017,-16'h0016,16'h001e,16'h001a,-16'h006e,16'h007d,16'h000e,-16'h002a,-16'h0013,16'h000d,-16'h0035,-16'h005e,16'h0017,-16'h000e,-16'h003f,16'h001d,16'h0081,-16'h0064,16'h002e,16'h0017,16'h0026,16'h002d,-16'h0019,-16'h0088,16'h003f,16'h0080,-16'h0002,16'h001c,16'h000c,16'h0039,-16'h0040,-16'h000e,16'h00a1,16'h0023,-16'h0015,16'h0058,16'h0003,-16'h000c,16'h000d,16'h0022,-16'h0040,-16'h001b,-16'h0006,-16'h001f,-16'h000d,16'h0018,16'h0049,16'h0044,16'h001e,16'h0035,-16'h0026,16'h0082,16'h002d,16'h0040,-16'h001e,-16'h0030,16'h003d,-16'h0030,16'h0029,-16'h0063,-16'h0032,-16'h002e,-16'h0035,16'h0016,16'h005e,-16'h004f,16'h004b,-16'h0036,16'h0009,-16'h0039,16'h0017,-16'h0031,-16'h002c,16'h000f,-16'h0046,-16'h0036,16'h0054,-16'h0021,-16'h001d,16'h000f,16'h0068,-16'h0088,16'h0042,16'h0017,-16'h0023,16'h004e,16'h0029,-16'h008a,16'h002c,16'h0044,16'h0048,16'h000f,-16'h001e,16'h001d,-16'h0041,-16'h002b,16'h00bc,16'h0032,-16'h0009,16'h003c,16'h0009,-16'h000d,16'h001a,16'h0023,-16'h004e,-16'h0031,16'h0019,-16'h0004,-16'h0045,16'h001c,16'h0039,16'h0027,16'h004c,16'h002f,-16'h0031,16'h0061,16'h0018,16'h0041,-16'h002f,-16'h0009,16'h003f,-16'h000f,16'h0023,-16'h00a7,-16'h005b,-16'h0026,16'h0003,16'h0001,16'h0047,-16'h002b,16'h0049,16'h0015,16'h0009,-16'h0026,16'h0004,-16'h0049,-16'h0029,16'h0021,-16'h006b,-16'h0032,16'h0061,-16'h0032,-16'h0029,16'h000d,16'h0054,-16'h00a3,16'h0037,16'h003e,-16'h0068,16'h0041,16'h000a,-16'h0021,16'h0046,16'h0035,16'h002b,-16'h0006,-16'h0035,16'h004f,-16'h002f,-16'h0033,16'h009f,16'h0045,-16'h001b,16'h005c,16'h0002,-16'h001f,-16'h002e,16'h0038,-16'h0026,-16'h0021,-16'h0002,16'h0006,-16'h0064,-16'h001a,16'h005f,16'h002c,16'h0070,16'h001f,-16'h0065,16'h0031,16'h0014,16'h0055,-16'h0033,-16'h0009,16'h0036,-16'h0033,16'h0061,-16'h00a8,-16'h008b,-16'h0016,-16'h0008,16'h000c,16'h004a,16'h0003,16'h0044,16'h0017,16'h000b,-16'h0013,16'h000b,-16'h003b,-16'h001d,16'h0057,-16'h00ab,-16'h001f,16'h0065,-16'h0037,-16'h0015,16'h0027,16'h002d,-16'h0078,16'h0018,16'h0041,-16'h00b1,16'h004a,16'h0005,16'h002e,16'h0035,16'h0002,16'h0045,-16'h000b,-16'h0040,16'h0056,-16'h0035,-16'h003e,16'h002d,16'h0011,-16'h0003,16'h005c,16'h000d,-16'h0012,-16'h002d,-16'h0008,-16'h0014,-16'h0024,-16'h000f,-16'h0009,-16'h0056,-16'h0012,16'h0076,16'h000c,16'h007a,16'h0044,-16'h003d,16'h002b,16'h0024,16'h0021,-16'h0084,-16'h000b,16'h003a,-16'h0035,16'h008e,-16'h008d,-16'h005b,-16'h001a,16'h0001,-16'h0024,16'h0060,16'h0013,16'h0061,16'h0049,16'h002c,16'h0005,16'h0016,-16'h002e,-16'h0055,16'h0051,-16'h00da,16'h0011,16'h004b,-16'h003d,-16'h0005,16'h003c,16'h001e,-16'h004b,-16'h000d,16'h0034,-16'h008c,16'h0063,16'h0008,16'h004f,16'h0021,-16'h0019,16'h0043,-16'h002c,-16'h0025,16'h0044,-16'h0025,-16'h002e,-16'h001f,16'h000a,-16'h0007,16'h0052,-16'h000f,16'h0007,-16'h000e,16'h0009,16'h0027,-16'h0022,-16'h0001,-16'h0028,-16'h0054,16'h0019,16'h0096,16'h0014,16'h007a,16'h0049,-16'h001e,16'h0038,16'h002b,16'h0023,-16'h0062,16'h000e,16'h0017,-16'h007a,16'h008b,-16'h006a,-16'h0039,16'h0004,16'h0024,-16'h0019,16'h0045,16'h003b,16'h004f,16'h0057,-16'h000c,-16'h0006,16'h0014,-16'h0031,-16'h0015,16'h0070,-16'h00b3,16'h0033,16'h0071,-16'h002f,-16'h0005,16'h0058,16'h0012,-16'h0010,16'h000c,16'h0000,-16'h00ac,16'h006b,-16'h0007,16'h0011,16'h0017,-16'h0015,16'h0050,-16'h0004,-16'h001f,16'h0055,16'h000e,-16'h0047,-16'h009d,16'h0014,16'h0000,16'h0056,-16'h0019,-16'h0003,-16'h0016,16'h0005,16'h0054,-16'h0009,16'h0008,-16'h0028,-16'h000d,16'h000f,16'h00a1,-16'h000f,16'h00a6,16'h004a,16'h0044,16'h0040,16'h0032,16'h003c,-16'h0081,16'h001f,-16'h000a,-16'h009f,16'h006f,-16'h0036,16'h0001,16'h002b,16'h0018,-16'h0031,16'h0030,16'h0031,16'h0039,16'h002a,-16'h0004,-16'h0005,16'h0017,-16'h0006,-16'h000d,16'h0085,-16'h0064,16'h003e,16'h0060,-16'h0021,-16'h001f,16'h001c,-16'h0008,16'h0006,16'h0013,16'h000d,-16'h0080,16'h0054,-16'h001a,-16'h0006,16'h0012,-16'h0035,16'h0068,-16'h0016,-16'h000c,16'h002b,-16'h0012,-16'h0030,-16'h0106,16'h004a,16'h0019,16'h0046,-16'h0015,16'h0005,-16'h0014,-16'h0007,16'h006e,-16'h0006,-16'h000b,-16'h0027,16'h0037,-16'h0002,16'h00b2,16'h0005,16'h00a8,16'h002b,16'h002f,16'h003a,16'h0034,16'h001e,-16'h006a,16'h001e,-16'h0038,-16'h00d1,16'h002c,-16'h001a,16'h0004,16'h0027,16'h0028,-16'h0027,-16'h0004,16'h0050,16'h003d,16'h0050,-16'h0016,-16'h000c,16'h002b,16'h0016,-16'h0016,16'h006b,16'h0006,16'h0001,16'h0041,-16'h0022,-16'h000d,16'h0011,-16'h0011,16'h0037,-16'h0010,-16'h0009,-16'h007a,16'h0028,-16'h0020,-16'h0042,16'h0010,-16'h0022,16'h0061,-16'h003e,16'h0006,16'h0012,-16'h002b,-16'h0076,-16'h011b,16'h003f,16'h0019,16'h001b,16'h0001,-16'h0020,-16'h002f,-16'h0001,16'h005f,-16'h0002,-16'h0006,-16'h0022,16'h005c,-16'h002a,16'h00c8,-16'h001e,16'h00a6,16'h003b,16'h0041,16'h002e,16'h0031,16'h0005,-16'h008f,16'h0016,-16'h001f,-16'h00d2,-16'h0022,16'h0012,-16'h0010,16'h0007,16'h0023,-16'h0022,-16'h000d,16'h0055,16'h0025,16'h0049,-16'h0012,-16'h0020,16'h000e,16'h000a,-16'h001a,16'h0054,16'h0034,16'h0007,16'h0040,-16'h0023,-16'h000e,16'h000a,-16'h0015,16'h0055,16'h000d,-16'h0010,-16'h0084,-16'h0008,-16'h001b,-16'h0062,-16'h0004,-16'h0043,16'h0058,-16'h0038,16'h0003,16'h0030,16'h0003,-16'h0089,-16'h00fd,16'h001a,-16'h0001,16'h0017,-16'h0023,-16'h0009,-16'h002d,-16'h0002,16'h0026,-16'h0022,-16'h0014,-16'h0005,16'h004f,-16'h0012,16'h00b7,-16'h0022,16'h009d,16'h0036,16'h002b,16'h0040,16'h003f,16'h0019,-16'h00d1,16'h0026,16'h0017,-16'h00aa,-16'h0059,16'h001d,-16'h0016,-16'h0025,16'h003d,-16'h001f,-16'h0029,16'h0019,16'h001e,16'h0049,-16'h0035,-16'h000c,16'h0000,16'h0003,-16'h0034,16'h0008,16'h0057,16'h000f,16'h0003,-16'h002c,16'h000d,-16'h0018,-16'h000e,16'h0059,16'h000a,-16'h003f,-16'h003d,-16'h0001,-16'h0015,-16'h003b,16'h0020,-16'h004a,16'h001b,-16'h0007,-16'h0006,16'h0048,16'h0021,-16'h009e,-16'h008f,16'h0030,16'h0005,16'h001b,-16'h0043,-16'h0010,-16'h0030,-16'h000c,16'h0061,-16'h0038,-16'h0009,16'h0005,16'h0076,16'h0012,16'h00c6,16'h0005,16'h0099,16'h002c,-16'h0005,16'h0043,16'h004b,16'h0004,-16'h017e,16'h0000,16'h0018,-16'h00c1,-16'h007d,16'h0015,-16'h0020,-16'h0034,16'h0029,16'h0000,-16'h0042,-16'h0013,16'h0033,16'h0039,-16'h000e,-16'h0010,16'h0003,-16'h000f,-16'h0015,16'h0003,16'h004d,-16'h002f,-16'h000b,-16'h001e,16'h0019,-16'h0009,-16'h0002,16'h0061,16'h001f,-16'h0032,-16'h002f,-16'h000c,-16'h001b,-16'h0017,-16'h0014,-16'h0035,16'h001a,-16'h0008,16'h0007,16'h003b,16'h0037,-16'h009f,-16'h0026,16'h002a,-16'h0009,16'h000a,-16'h001a,-16'h0006,-16'h0027,-16'h0014,16'h005a,-16'h0037,-16'h0032,16'h0022,16'h0047,16'h0024,16'h00c1,-16'h0024,16'h00a9,16'h004b,16'h0016,16'h0045,16'h002c,-16'h0022,-16'h014d,16'h0020,-16'h0011,-16'h0092,-16'h0059,16'h0011,-16'h0027,-16'h002b,16'h0035,16'h0009,-16'h0011,-16'h0072,16'h003f,16'h0021,-16'h0017,-16'h0021,-16'h0001,16'h0012,-16'h0018,-16'h0018,16'h003f,-16'h0022,-16'h001d,-16'h0010,16'h003f,16'h0000,-16'h0005,16'h0079,16'h0008,-16'h0033,-16'h001f,-16'h000b,-16'h000a,16'h0064,-16'h0010,-16'h0014,16'h0002,-16'h0017,-16'h0018,16'h0036,16'h0050,-16'h0060,16'h001e,16'h0012,-16'h0021,16'h001f,-16'h0002,-16'h0010,-16'h0039,-16'h001e,16'h004a,-16'h0027,-16'h001c,16'h0031,-16'h0005,16'h0008,16'h00a7,-16'h004c,16'h0099,16'h003d,16'h0011,16'h002b,16'h004e,-16'h000d,-16'h00ef,16'h0005,16'h0017,-16'h0082,-16'h0055,-16'h0015,-16'h0017,-16'h0033,16'h003a,16'h0005,-16'h0028,-16'h0055,16'h0042,16'h0012,-16'h0010,-16'h0010,-16'h0003,-16'h0021,16'h0004,-16'h0034,16'h0049,-16'h0014,-16'h000e,16'h0002,16'h0017,-16'h0008,16'h0006,16'h0076,-16'h000f,-16'h0010,-16'h0018,-16'h002c,-16'h0021,16'h0065,-16'h0018,-16'h0020,16'h0007,-16'h0012,-16'h000b,16'h002b,16'h005b,-16'h0022,16'h003e,-16'h001b,-16'h0022,16'h0020,-16'h0009,-16'h0005,16'h0018,-16'h001a,16'h004d,-16'h0026,-16'h0020,16'h0003,-16'h002f,-16'h000f,16'h00ab,-16'h0008,16'h0088,16'h0051,16'h0028,16'h0004,16'h0042,16'h0003,-16'h005a,-16'h000f,16'h001e,-16'h008f,-16'h005a,-16'h0005,-16'h0010,-16'h004d,16'h0000,16'h002c,-16'h0029,-16'h004a,16'h0052,16'h0011,-16'h0010,-16'h0022,16'h0004,-16'h0020,16'h001c,-16'h001f,16'h0033,-16'h0013,16'h000f,-16'h0002,16'h000b,-16'h0021,16'h0003,16'h008c,-16'h0009,16'h000a,-16'h003b,-16'h0031,16'h0007,16'h006f,16'h002e,16'h000d,-16'h0003,-16'h000c,-16'h0013,16'h0024,16'h005a,16'h0013,16'h004b,16'h001b,-16'h001c,16'h002a,16'h0018,-16'h0006,16'h003a,-16'h001a,16'h0030,-16'h0053,-16'h0032,-16'h001e,-16'h0036,-16'h0019,16'h009c,16'h002a,16'h0086,16'h006b,16'h0011,16'h0007,16'h0032,-16'h000a,-16'h0052,-16'h0014,16'h003a,-16'h0095,-16'h005b,-16'h0015,16'h0026,-16'h003c,16'h0037,16'h003c,-16'h0011,-16'h0019,16'h005d,-16'h0029,16'h0001,-16'h0010,16'h0000,-16'h003e,-16'h000a,-16'h0015,16'h0036,16'h0018,16'h0016,16'h001c,16'h0000,-16'h001a,-16'h0003,16'h0088,16'h0011,16'h0006,-16'h0020,-16'h0046,16'h0026,16'h001e,16'h0040,16'h0030,16'h0022,-16'h000b,-16'h0018,16'h001d,16'h005a,16'h0057,16'h004a,16'h002b,-16'h0004,16'h000e,-16'h0004,-16'h0002,16'h0011,-16'h0013,16'h0036,-16'h0042,-16'h0024,-16'h0012,-16'h0036,-16'h001e,16'h0083,16'h0038,16'h0094,16'h00a2,16'h001c,-16'h0015,16'h002a,16'h000b,-16'h0056,-16'h0006,16'h003f,-16'h0076,-16'h0058,16'h0019,16'h0011,-16'h004d,16'h0036,16'h0033,-16'h0012,16'h0029,16'h0055,-16'h0033,-16'h0001,-16'h003f,-16'h0001,-16'h0025,16'h0000,16'h0005,16'h0047,16'h0013,-16'h000a,16'h0000,16'h0010,-16'h000c,-16'h000d,16'h005d,16'h0000,16'h0019,16'h003e,-16'h0021,16'h0003,-16'h006d,16'h0052,16'h002a,16'h000d,-16'h0003,-16'h000f,16'h001b,16'h0036,16'h0042,16'h0057,16'h0026,16'h000c,16'h0016,-16'h0002,-16'h0005,-16'h0028,-16'h000c,16'h003b,-16'h0011,-16'h0020,-16'h000a,-16'h0010,-16'h0038,16'h007b,16'h0036,16'h0068,16'h0094,16'h000d,-16'h0015,16'h003a,16'h001d,-16'h006e,-16'h000d,16'h003b,-16'h007b,-16'h005f,16'h0016,-16'h000c,-16'h0073,16'h001a,16'h0022,16'h000c,16'h0046,16'h0043,-16'h0011,16'h0005,-16'h001d,-16'h0007,-16'h0007,-16'h000b,16'h0002,16'h006e,16'h002f,16'h0004,-16'h0005,16'h0019,-16'h0008,-16'h0018,16'h0012,-16'h0004,16'h0042,16'h004c,-16'h0036,16'h0028,-16'h009e,16'h0061,16'h005f,16'h000f,16'h0005,-16'h0010,16'h0025,-16'h001d,16'h005c,16'h0039,16'h0025,-16'h0018,16'h001d,16'h0001,16'h0001,-16'h0057,16'h0001,16'h0035,16'h001e,-16'h002c,16'h0022,-16'h0009,-16'h0009,16'h007b,16'h003d,16'h0070,16'h0093,-16'h0009,-16'h0026,-16'h000e,16'h0048,-16'h0047,-16'h004a,16'h0038,-16'h006b,-16'h0037,16'h002d,-16'h0017,-16'h007c,16'h0035,16'h0042,16'h0004,16'h003b,16'h0060,-16'h002b,16'h0021,-16'h0023,-16'h0007,-16'h0007,-16'h000a,-16'h0008,16'h0083,16'h004b,-16'h0034,-16'h0014,16'h0037,-16'h0017,16'h0005,-16'h001a,-16'h001e,16'h0030,16'h004a,-16'h001d,16'h000d,-16'h005c,16'h0070,16'h007f,16'h0022,16'h000d,-16'h000b,16'h003d,-16'h00ab,16'h0063,16'h0017,-16'h0016,-16'h0015,-16'h0017,-16'h0008,-16'h0012,-16'h006d,-16'h0007,-16'h0011,16'h0024,-16'h002f,16'h0041,16'h0015,16'h0030,16'h0072,16'h004f,16'h004c,16'h0067,16'h0007,-16'h003c,-16'h0011,16'h0029,16'h0001,-16'h0027,16'h0037,-16'h005f,-16'h0047,16'h0036,-16'h0025,-16'h0056,16'h0052,16'h0066,-16'h0014,16'h0026,16'h004f,-16'h0023,16'h005d,-16'h002c,16'h0009,16'h0002,-16'h000b,16'h000b,16'h0059,16'h005d,-16'h0034,-16'h000e,16'h0014,-16'h005d,16'h0005,-16'h0053,-16'h001c,16'h001e,16'h0053,16'h002c,-16'h0004,-16'h0025,16'h0057,16'h008a,-16'h0003,16'h0001,-16'h000d,16'h0066,-16'h0187,16'h0059,16'h0002,-16'h000f,-16'h0008,-16'h0005,-16'h000a,-16'h0027,-16'h003d,-16'h0009,-16'h0026,16'h0027,16'h000b,16'h004f,-16'h0028,16'h0062,16'h0074,-16'h001b,16'h0062,16'h0055,16'h0000,-16'h0026,-16'h0001,-16'h0057,16'h0058,-16'h0046,16'h002f,-16'h0062,-16'h0052,16'h0046,-16'h000f,-16'h0043,16'h0050,16'h006a,16'h0008,16'h0036,16'h005f,-16'h0014,16'h0058,-16'h0014,16'h000c,-16'h0007,16'h0019,16'h000e,16'h0075,16'h0053,-16'h0028,-16'h0012,16'h002a,-16'h0054,16'h0006,-16'h006d,-16'h0002,16'h0029,16'h0063,16'h0048,16'h0019,-16'h000e,16'h0038,16'h0081,-16'h0037,16'h0011,-16'h000d,16'h0060,-16'h01fe,16'h0028,-16'h000e,-16'h000d,-16'h000b,16'h0004,-16'h000f,-16'h0032,16'h001a,16'h000b,-16'h0040,16'h0001,16'h0030,16'h002e,-16'h0030,16'h0057,16'h0091,-16'h0088,16'h0069,16'h0057,-16'h000d,-16'h0009,-16'h0012,-16'h0121,16'h004d,-16'h0036,16'h0034,-16'h0066,-16'h0057,16'h002d,-16'h0002,-16'h0038,16'h0025,16'h0073,16'h0038,16'h0023,16'h005d,-16'h001e,16'h0052,16'h0007,16'h0007,16'h0009,16'h0020,-16'h0020,16'h0091,16'h004e,-16'h004b,-16'h0021,16'h0039,-16'h002d,-16'h0013,-16'h00a9,-16'h001d,16'h0022,16'h006b,16'h0056,16'h000c,16'h0027,-16'h002b,16'h006c,-16'h007f,16'h0011,-16'h0001,16'h004a,-16'h017c,-16'h0011,-16'h001f,16'h0035,-16'h0008,-16'h000d,16'h0011,-16'h0044,16'h006d,16'h0020,-16'h005c,16'h001c,16'h001b,16'h0048,-16'h0034,16'h0037,16'h0052,-16'h0088,16'h003b,16'h0042,16'h0007,16'h003b,-16'h0001,-16'h0179,16'h006e,-16'h007c,16'h0037,-16'h0069,-16'h0044,16'h0011,16'h0011,-16'h0036,16'h0033,16'h005e,16'h0042,16'h0026,16'h0058,16'h0013,16'h0048,16'h000f,16'h0024,-16'h0024,16'h002b,16'h0000,16'h009d,16'h0041,-16'h005a,-16'h0020,16'h003b,-16'h003d,-16'h0013,-16'h00ac,16'h0004,16'h001e,16'h0038,16'h002c,16'h0014,16'h0005,-16'h00b7,16'h0056,-16'h006f,-16'h000f,16'h0030,16'h001e,-16'h00b5,-16'h001e,-16'h0022,16'h0034,-16'h0019,16'h0008,16'h005c,-16'h002c,16'h0081,-16'h000e,-16'h00a5,16'h0007,16'h0000,16'h001e,-16'h002a,-16'h0017,16'h0026,-16'h0009,16'h005d,16'h0046,16'h0007,16'h0058,-16'h0021,-16'h0162,16'h0047,-16'h008b,16'h000a,-16'h005f,-16'h000b,16'h0028,-16'h0004,-16'h0027,16'h004d,16'h0055,16'h002c,-16'h0002,16'h0049,16'h0009,16'h002f,16'h000c,16'h001b,-16'h000f,16'h0052,-16'h0009,16'h0072,16'h003d,-16'h002f,-16'h0014,16'h002a,-16'h000e,16'h0014,-16'h00cf,16'h0015,16'h001f,16'h0018,16'h0033,16'h0049,-16'h001c,-16'h0103,16'h0058,-16'h0054,-16'h0008,16'h000d,16'h0037,-16'h0077,-16'h000f,-16'h000d,16'h0047,16'h000d,-16'h0002,16'h0077,-16'h0041,16'h0021,-16'h000d,-16'h00b3,16'h0001,-16'h001f,16'h0026,16'h000a,-16'h004c,16'h0048,16'h005b,16'h004b,16'h0047,16'h0025,16'h0067,-16'h0019,-16'h012d,16'h0055,-16'h0088,-16'h0005,-16'h005f,16'h0038,16'h0023,16'h0000,-16'h0035,16'h0043,16'h003f,16'h0015,-16'h001b,16'h005f,-16'h0003,16'h0034,16'h0041,16'h0016,16'h000a,16'h0047,16'h0012,16'h008f,16'h0054,-16'h0012,16'h0006,16'h002f,16'h0003,-16'h0016,-16'h00d8,16'h0024,16'h0020,-16'h001b,16'h003f,16'h0034,-16'h0007,-16'h00c3,16'h005d,-16'h000c,16'h0000,16'h001a,16'h0030,-16'h004b,-16'h0015,-16'h0033,16'h002b,-16'h0005,-16'h0009,16'h006b,-16'h0048,-16'h0011,-16'h001d,-16'h00ae,-16'h001c,-16'h005b,16'h005c,16'h000f,-16'h0052,16'h0045,16'h00c5,16'h003a,16'h0047,16'h002d,16'h0057,-16'h0010,-16'h00e3,16'h0042,-16'h0046,-16'h0022,-16'h004d,16'h003b,16'h0016,-16'h000b,-16'h0009,16'h003c,16'h0038,16'h002f,-16'h0013,16'h0085,-16'h0013,16'h0054,16'h0051,16'h0014,16'h0000,16'h0049,16'h001a,16'h006b,16'h004d,16'h0003,16'h0024,16'h0036,16'h0004,16'h0008,-16'h00dc,16'h001c,16'h001e,-16'h006b,16'h004f,16'h0033,16'h0016,-16'h0050,16'h0077,16'h000e,16'h0007,16'h0004,16'h003f,-16'h0034,16'h000a,-16'h002d,16'h0001,-16'h002e,-16'h0017,16'h0034,-16'h003a,-16'h0035,-16'h0036,-16'h007c,-16'h0003,-16'h00ad,16'h0021,-16'h0027,-16'h0039,16'h0062,16'h00e7,16'h0041,16'h0053,16'h0036,16'h0072,-16'h0002,-16'h0075,16'h0044,-16'h001c,-16'h0042,-16'h002b,16'h0034,16'h0044,16'h0001,16'h0010,16'h0025,-16'h0065,16'h0055,-16'h0021,16'h009e,16'h000d,16'h006e,16'h0045,-16'h0021,-16'h0013,16'h003c,16'h003b,16'h002d,16'h0046,16'h0001,16'h0036,16'h003d,16'h0047,16'h000f,-16'h00d3,-16'h0008,16'h0031,-16'h00dd,16'h0059,16'h0026,-16'h0021,16'h0017,16'h0080,16'h005e,16'h0011,-16'h000a,16'h001b,-16'h001e,-16'h0014,-16'h003f,-16'h002e,-16'h0031,-16'h0013,16'h002f,-16'h0059,-16'h0075,-16'h0034,-16'h0039,-16'h0012,-16'h00a1,16'h0021,-16'h0022,-16'h0003,16'h0071,16'h00a7,16'h004c,16'h004d,16'h0040,16'h005b,16'h0002,-16'h0048,16'h002a,-16'h0015,-16'h002f,-16'h001b,16'h002d,16'h005d,-16'h0009,16'h0022,-16'h0016,-16'h00a3,16'h0053,-16'h0011,16'h0076,16'h001f,16'h004c,16'h0074,-16'h0029,-16'h0030,16'h002b,16'h0029,16'h000f,16'h0020,-16'h000f,16'h001d,16'h002f,16'h0046,16'h0037,-16'h0092,16'h0029,16'h0040,-16'h0132,16'h007a,16'h001e,-16'h001a,16'h0068,16'h0077,16'h0075,-16'h0011,-16'h003b,16'h0027,-16'h0014,-16'h0036,-16'h0025,-16'h0042,-16'h0012,16'h0013,16'h0023,-16'h002c,-16'h008b,16'h0040,-16'h0022,16'h0015,-16'h00b7,16'h0023,-16'h001b,-16'h0013,16'h00b9,16'h004c,16'h0015,16'h002a,16'h0040,16'h0073,16'h000f,-16'h004e,16'h0055,16'h0015,16'h0003,-16'h0022,16'h002f,16'h0067,-16'h001e,-16'h0021,-16'h0053,-16'h00cb,16'h0051,-16'h000d,16'h0040,16'h0011,-16'h0029,16'h0079,-16'h001a,-16'h001e,-16'h0009,16'h0020,-16'h0006,16'h0046,-16'h000d,16'h0033,16'h002e,16'h0054,16'h0015,-16'h0083,16'h0023,16'h002a,-16'h010b,16'h0033,16'h0014,16'h0010,16'h0077,16'h006e,16'h0071,16'h001f,-16'h0039,16'h0022,-16'h0009,-16'h0046,-16'h0047,-16'h002f,-16'h0010,16'h0022,16'h0028,-16'h0018,-16'h0050,16'h002d,-16'h0028,-16'h0004,-16'h0080,16'h0029,-16'h0014,-16'h0016,16'h00b5,16'h001f,16'h0010,16'h001f,16'h0076,16'h0075,16'h003a,-16'h003b,16'h004a,16'h0048,-16'h0013,-16'h0010,16'h0051,16'h007c,-16'h0037,-16'h0007,-16'h0030,-16'h0085,16'h0044,16'h0010,16'h0038,16'h0007,-16'h006b,16'h007c,16'h000e,-16'h000e,-16'h0008,-16'h0004,-16'h0042,-16'h0086,16'h0000,-16'h0007,16'h0004,16'h001d,16'h00a7,-16'h0055,16'h0036,16'h000f,16'h001a,16'h0033,16'h0005,-16'h0081,16'h0038,16'h0072,-16'h0006,-16'h0017,-16'h0005,16'h004a,-16'h0048,16'h0000,16'h00bb,16'h0057,-16'h002a,16'h004a,16'h002b,-16'h002e,16'h002e,16'h002e,-16'h0037,-16'h0017,16'h0013,-16'h0002,-16'h0027,16'h001f,16'h0021,16'h006c,16'h004f,16'h002c,-16'h002f,16'h0057,16'h0010,16'h006d,-16'h004b,-16'h0032,16'h0047,-16'h0007,16'h0019,-16'h007d,-16'h002f,-16'h0044,-16'h001a,-16'h0006,16'h0053,-16'h0027,16'h0038,16'h0003,16'h0027,-16'h002f,16'h0023,-16'h0037,-16'h0008,16'h002e,-16'h0054,-16'h0047,16'h0000,-16'h0026,16'h001b,16'h000e,16'h0087,-16'h008c,16'h0055,16'h0032,-16'h0016,16'h001b,16'h0018,-16'h0042,16'h0029,16'h0048,16'h0001,-16'h000d,-16'h002f,16'h0031,-16'h0036,-16'h001b,16'h00ab,16'h0039,16'h000b,16'h0073,16'h0001,-16'h001d,16'h000d,16'h0004,-16'h003d,-16'h001f,16'h001f,-16'h0013,-16'h0035,16'h0010,16'h0014,16'h0031,16'h0061,16'h002c,-16'h0059,16'h0041,16'h0005,16'h005b,-16'h004a,-16'h000f,16'h0053,-16'h002e,16'h0056,-16'h008f,-16'h005d,-16'h002e,-16'h0006,16'h000e,16'h0045,16'h000d,16'h0034,16'h000a,16'h000c,-16'h0015,16'h001a,-16'h0024,-16'h0027,16'h0042,-16'h0080,-16'h002a,16'h0008,-16'h0041,16'h000c,16'h0012,16'h0049,-16'h008f,16'h002c,16'h006a,-16'h005f,16'h0054,-16'h000a,16'h001b,16'h001b,16'h0022,-16'h0004,-16'h001d,-16'h001b,16'h0020,-16'h0042,-16'h000c,16'h006f,16'h0032,-16'h001d,16'h008d,16'h0008,-16'h0040,-16'h0029,16'h0023,-16'h001e,-16'h001b,16'h0018,-16'h0012,-16'h0039,-16'h002f,16'h0009,16'h0029,16'h0099,16'h0017,-16'h0069,16'h002b,16'h0009,16'h0048,-16'h007b,16'h000e,16'h0038,-16'h0019,16'h0080,-16'h0062,-16'h0037,-16'h002c,16'h002d,-16'h001a,16'h0038,16'h0019,16'h0043,16'h000a,-16'h001b,-16'h0021,16'h0026,-16'h002b,-16'h0045,16'h006b,-16'h00a8,-16'h0002,16'h0014,-16'h0029,-16'h000d,16'h0038,16'h0024,-16'h0061,16'h000c,16'h004c,-16'h005d,16'h0034,16'h0013,16'h0040,16'h0001,16'h0018,16'h000e,-16'h000a,-16'h0037,16'h004a,-16'h0017,-16'h0012,16'h002f,16'h0014,-16'h0004,16'h008c,-16'h0013,-16'h000a,-16'h002e,-16'h0003,16'h001c,-16'h0013,16'h000e,-16'h0023,-16'h0030,-16'h0019,16'h004d,16'h0007,16'h0089,16'h0030,-16'h005c,16'h002c,16'h0017,16'h0040,-16'h007c,16'h0004,16'h0029,-16'h0036,16'h0098,-16'h0043,-16'h0046,16'h0009,-16'h0003,16'h0000,16'h004d,16'h0030,16'h001a,16'h0040,16'h000b,-16'h0012,16'h0047,-16'h0045,-16'h004b,16'h0078,-16'h00cb,16'h0028,-16'h0003,-16'h0012,16'h0002,16'h0026,16'h0009,-16'h003c,-16'h0023,16'h0032,-16'h007d,16'h0058,-16'h001a,16'h0037,-16'h002d,16'h0007,16'h0020,-16'h0007,-16'h0030,16'h003d,-16'h0005,-16'h0024,-16'h003a,16'h0011,-16'h0026,16'h0042,-16'h002a,16'h000e,-16'h0021,16'h0002,16'h0043,-16'h0011,-16'h0010,-16'h002f,-16'h003e,16'h0012,16'h0075,16'h0003,16'h00a2,16'h0044,-16'h001b,16'h0048,16'h002f,16'h0038,-16'h0078,16'h001a,16'h0031,-16'h0055,16'h009a,-16'h000d,-16'h0027,16'h003d,16'h0019,16'h0001,16'h0026,16'h0056,16'h002e,16'h003b,-16'h000d,-16'h0011,16'h005b,-16'h0027,-16'h003d,16'h006f,-16'h0073,16'h0024,-16'h002c,-16'h003a,16'h000b,16'h0033,16'h0000,-16'h0017,16'h0004,16'h0018,-16'h0058,16'h0035,-16'h000d,16'h000e,-16'h001d,16'h0006,16'h0006,-16'h0020,-16'h0012,16'h0034,-16'h0016,-16'h0040,-16'h00a8,16'h0032,16'h000d,16'h0062,-16'h000c,16'h0012,-16'h0001,-16'h000a,16'h0060,16'h0015,16'h002f,-16'h0041,16'h0010,16'h0008,16'h0089,16'h000c,16'h00aa,16'h0035,16'h0017,16'h0023,16'h000d,16'h0035,-16'h008e,16'h002e,16'h0007,-16'h006b,16'h006d,-16'h0018,-16'h001c,16'h004c,16'h0023,-16'h0028,16'h0015,16'h0031,16'h0033,16'h0036,-16'h0006,-16'h0009,16'h004c,-16'h0036,-16'h002a,16'h007f,-16'h001a,16'h0009,-16'h0047,-16'h003b,16'h0013,16'h0036,-16'h0006,16'h0033,-16'h000d,16'h0005,-16'h005f,16'h002a,-16'h0025,-16'h0030,-16'h001c,-16'h0019,16'h000b,-16'h0053,-16'h0023,16'h0027,-16'h0041,-16'h0053,-16'h0110,16'h0046,-16'h0010,16'h003e,16'h0002,-16'h0008,-16'h0012,-16'h000b,16'h0048,-16'h000a,16'h0027,-16'h002f,16'h0049,-16'h0009,16'h0093,16'h0000,16'h00bf,16'h0025,16'h0029,16'h0033,16'h0029,16'h0047,-16'h009d,16'h0025,-16'h000a,-16'h008f,16'h0039,-16'h000a,-16'h0013,16'h0033,16'h0016,-16'h002a,-16'h000b,16'h0061,16'h0032,16'h005a,-16'h001b,-16'h0027,16'h0052,-16'h0009,-16'h0032,16'h0045,16'h0028,16'h000b,-16'h003e,-16'h002b,16'h0007,16'h0019,16'h0007,16'h007a,-16'h0016,16'h000f,-16'h0079,16'h0027,-16'h003f,-16'h007b,-16'h0012,-16'h0013,16'h0020,-16'h002f,-16'h0005,16'h0048,-16'h0036,-16'h0048,-16'h013c,16'h003f,-16'h001e,16'h0054,-16'h0009,-16'h0008,-16'h0015,-16'h0026,16'h004c,16'h000a,-16'h000b,-16'h0019,16'h0025,-16'h0013,16'h00aa,16'h0000,16'h00ab,16'h0007,16'h002e,16'h0045,16'h0023,16'h003a,-16'h00de,16'h0008,16'h0014,-16'h0086,-16'h0030,-16'h0012,-16'h003f,16'h004c,16'h0025,-16'h000b,-16'h0033,16'h0021,16'h002e,16'h003d,-16'h0015,-16'h0027,16'h0041,-16'h0012,-16'h0036,16'h0024,16'h006c,-16'h000f,-16'h008f,-16'h0022,-16'h0018,-16'h0014,-16'h000a,16'h0080,-16'h0028,16'h000e,-16'h0068,16'h001b,-16'h0028,-16'h0081,16'h0002,-16'h0011,16'h003d,-16'h0020,16'h0007,16'h001a,-16'h001b,-16'h009d,-16'h00ad,16'h0047,16'h0003,16'h003c,-16'h0015,-16'h0001,-16'h002b,-16'h0018,16'h0054,-16'h0032,16'h0002,-16'h000c,16'h0033,16'h0017,16'h00ab,-16'h0027,16'h00ab,16'h0000,16'h0029,16'h0033,16'h0003,16'h001a,-16'h0156,-16'h000b,16'h0009,-16'h0028,-16'h0054,16'h0006,-16'h0011,16'h002b,16'h0033,16'h000f,-16'h004b,-16'h003c,16'h0029,16'h002c,-16'h0035,-16'h0026,16'h0035,-16'h0005,-16'h001d,16'h0041,16'h0048,-16'h000e,-16'h0096,-16'h000a,-16'h0025,-16'h0005,-16'h0005,16'h00a8,-16'h0019,-16'h000e,-16'h002e,16'h0027,-16'h0017,-16'h0038,-16'h000c,-16'h001f,16'h0028,-16'h0007,16'h0004,16'h004e,16'h001e,-16'h00b9,-16'h002a,16'h003d,-16'h0003,16'h0020,16'h0002,-16'h001c,-16'h0060,-16'h0003,16'h006a,-16'h001c,-16'h0029,16'h0009,16'h0055,16'h0026,16'h00db,-16'h000f,16'h00b4,16'h000c,-16'h0009,16'h0053,16'h0028,-16'h0004,-16'h0160,16'h0003,16'h0024,-16'h001a,-16'h0070,-16'h001d,-16'h0009,16'h0019,16'h002e,16'h0003,-16'h0066,-16'h0075,16'h002d,16'h002f,-16'h002e,-16'h000e,16'h0012,16'h0003,-16'h002c,16'h000c,16'h0023,-16'h0035,-16'h0070,-16'h0018,-16'h0013,16'h0000,-16'h0014,16'h00ab,-16'h0009,16'h0000,-16'h0037,16'h0014,-16'h0031,16'h0039,-16'h002b,16'h0000,-16'h0009,-16'h0011,16'h0009,16'h0042,16'h0030,-16'h00b3,16'h0012,16'h0029,16'h0009,16'h0040,-16'h0004,-16'h0019,-16'h004f,-16'h000b,16'h006b,16'h0004,-16'h0042,16'h002b,16'h001f,16'h0001,16'h00d3,-16'h0023,16'h0093,16'h0047,16'h000f,16'h0044,16'h003b,16'h0022,-16'h010b,-16'h0008,16'h0005,-16'h0037,-16'h0076,-16'h000d,16'h0003,16'h002d,16'h0046,16'h000b,-16'h0049,-16'h0079,16'h0034,16'h0008,-16'h0029,-16'h002d,16'h0033,-16'h000c,-16'h001f,-16'h0023,16'h0028,-16'h0020,-16'h0086,16'h0001,-16'h001e,16'h0005,16'h000d,16'h007e,16'h0010,-16'h0029,-16'h001a,16'h0035,-16'h0025,16'h0086,-16'h004e,16'h0006,-16'h001c,16'h0005,-16'h0001,16'h003f,16'h0051,-16'h0053,16'h0023,-16'h0009,-16'h003c,16'h0032,16'h0018,-16'h0002,-16'h001d,16'h0016,16'h005d,-16'h0010,-16'h003f,16'h0013,-16'h0034,16'h000e,16'h00df,-16'h0045,16'h0099,16'h0034,16'h0024,16'h003d,16'h0030,16'h0027,-16'h00aa,-16'h0007,16'h0024,-16'h0031,-16'h007a,-16'h000e,-16'h0018,16'h0011,16'h0044,-16'h001c,-16'h0050,-16'h005b,16'h0059,16'h0013,-16'h0009,-16'h0024,16'h000a,-16'h001e,16'h0007,-16'h001c,16'h0031,-16'h0009,-16'h00a6,16'h0004,-16'h0005,-16'h000b,16'h0031,16'h0087,16'h000b,-16'h0010,-16'h002a,16'h000b,-16'h0011,16'h0080,-16'h0039,-16'h0004,-16'h0007,-16'h0006,16'h0010,16'h003d,16'h007b,-16'h0001,16'h0051,-16'h0011,-16'h0010,16'h0051,-16'h000c,-16'h0001,-16'h0009,16'h0007,16'h006d,-16'h002e,-16'h0030,16'h000e,-16'h0083,16'h0017,16'h00c9,16'h0000,16'h0092,16'h002c,16'h000b,16'h0015,16'h0025,16'h0009,-16'h0027,-16'h0021,16'h004a,-16'h0031,-16'h008b,-16'h0022,16'h0014,16'h0023,16'h0031,16'h0012,-16'h0042,-16'h0006,16'h007c,-16'h0010,16'h0009,-16'h000f,-16'h001a,-16'h0006,-16'h0016,-16'h0017,16'h002d,16'h0017,-16'h0089,16'h0013,16'h0008,16'h0000,16'h000c,16'h0072,-16'h0002,16'h0006,-16'h0039,-16'h002e,-16'h002c,16'h0049,16'h0012,16'h0031,-16'h001a,-16'h000e,16'h0002,16'h001f,16'h0086,16'h005e,16'h0029,16'h0017,-16'h0008,16'h0035,16'h0010,-16'h0024,16'h0028,-16'h000f,16'h0051,-16'h0035,-16'h0047,-16'h001b,-16'h0070,16'h0000,16'h00bb,16'h0017,16'h0098,16'h0038,16'h000d,16'h0027,16'h0033,16'h002f,-16'h0045,-16'h0005,16'h0020,-16'h004e,-16'h0091,-16'h0002,16'h0015,-16'h0002,16'h004a,16'h0022,-16'h0034,16'h0024,16'h0079,-16'h002c,16'h0019,16'h000c,16'h0002,-16'h002b,-16'h000e,-16'h000f,16'h0045,16'h0035,-16'h008a,-16'h0009,-16'h0017,16'h0011,16'h000c,16'h0046,16'h0006,16'h000e,-16'h002b,-16'h0036,16'h0003,-16'h0037,16'h0048,16'h005a,16'h0017,16'h0009,-16'h000a,16'h000f,16'h00ab,16'h0065,16'h0051,16'h001e,16'h0007,16'h0031,16'h000a,16'h0012,16'h000a,-16'h001d,16'h005d,-16'h0013,-16'h004a,-16'h003a,-16'h001f,-16'h0024,16'h0087,16'h002b,16'h0099,16'h0057,-16'h0006,16'h0015,16'h0040,16'h0014,-16'h005b,-16'h0018,16'h003a,-16'h0004,-16'h0063,16'h0020,16'h0018,-16'h0019,16'h0040,16'h0011,-16'h0018,16'h0055,16'h006a,-16'h002a,16'h0019,-16'h0006,16'h001f,-16'h001e,16'h0010,-16'h0007,16'h006f,16'h005e,-16'h007d,16'h0016,16'h0019,16'h0004,-16'h0002,-16'h0004,-16'h001b,16'h0015,16'h0030,-16'h0033,16'h0014,-16'h006a,16'h004e,16'h0049,16'h001c,-16'h0004,16'h0005,16'h000f,16'h006c,16'h0061,16'h0038,16'h0017,-16'h000b,16'h0042,16'h0011,-16'h000c,-16'h0023,-16'h0007,16'h002f,16'h0021,-16'h0021,16'h0001,-16'h0003,-16'h0049,16'h0076,16'h0049,16'h0095,16'h0065,16'h0011,16'h000d,16'h001d,16'h0045,-16'h003e,16'h0004,16'h0033,-16'h0007,-16'h0013,16'h0042,16'h0025,-16'h0019,16'h0042,16'h003d,-16'h003a,16'h005d,16'h006d,-16'h003e,16'h0012,-16'h000f,-16'h0007,-16'h0013,-16'h0003,16'h0013,16'h007a,16'h0063,-16'h00b0,16'h0018,16'h002c,-16'h000e,16'h0016,-16'h0015,16'h0009,16'h0024,16'h0063,-16'h0024,16'h0026,-16'h009e,16'h0084,16'h0066,-16'h0006,16'h0024,-16'h0002,16'h0026,16'h0016,16'h0044,16'h0027,16'h002f,-16'h0029,16'h0041,16'h001e,-16'h000f,-16'h0096,16'h0011,16'h000a,16'h002b,-16'h0027,16'h0018,16'h0018,-16'h0039,16'h006a,16'h003b,16'h0074,16'h005f,16'h0002,-16'h0021,16'h0023,16'h0065,-16'h0036,-16'h002f,16'h002e,16'h0027,-16'h0055,16'h004f,16'h001f,-16'h001c,16'h0046,16'h0054,-16'h004a,16'h0015,16'h005d,-16'h0024,16'h0006,-16'h0006,-16'h000b,-16'h000f,-16'h002c,16'h0009,16'h0072,16'h0061,-16'h00ae,16'h000f,16'h0017,16'h0005,16'h0007,-16'h005e,-16'h0027,16'h002e,16'h006b,-16'h001c,16'h0046,-16'h002e,16'h0091,16'h0099,-16'h000e,16'h002d,-16'h002c,16'h003e,-16'h008c,16'h0065,16'h001a,16'h0006,-16'h000e,16'h0026,16'h0012,-16'h0022,-16'h008e,-16'h0004,-16'h002b,16'h0014,-16'h0015,16'h0036,-16'h000d,16'h0014,16'h006e,16'h0038,16'h0068,16'h0041,-16'h0007,-16'h001b,16'h0009,16'h004c,16'h0021,-16'h0025,16'h0038,16'h0021,-16'h004b,16'h0060,16'h0002,-16'h003b,16'h0036,16'h004b,-16'h003d,16'h000c,16'h0053,16'h0000,16'h0049,-16'h0033,16'h0005,-16'h0013,-16'h0028,16'h000f,16'h0062,16'h005b,-16'h00a9,-16'h000a,16'h003b,-16'h002f,16'h0005,-16'h0082,-16'h0010,16'h0015,16'h0048,16'h0007,16'h0026,-16'h002b,16'h0078,16'h009c,-16'h000e,16'h0007,-16'h0008,16'h005c,-16'h01a3,16'h0029,-16'h0006,-16'h0004,-16'h0006,16'h0014,16'h000c,-16'h0020,-16'h0063,16'h0008,-16'h0041,16'h0021,16'h0004,16'h0033,-16'h003c,16'h0046,16'h0057,16'h0003,16'h0063,16'h0024,-16'h000c,-16'h0011,16'h002c,16'h0015,16'h003a,-16'h0019,16'h002c,16'h0002,-16'h006b,16'h0066,-16'h0004,-16'h0027,16'h0042,16'h0045,-16'h000f,16'h000b,16'h005a,16'h000f,16'h005b,-16'h0015,16'h000b,-16'h0016,16'h001b,16'h0007,16'h006c,16'h005e,-16'h0097,-16'h001d,16'h003b,-16'h0021,16'h001a,-16'h0096,-16'h000e,-16'h002b,16'h006b,16'h002d,16'h0014,16'h000c,16'h0035,16'h0099,-16'h0037,16'h000f,-16'h0019,16'h0058,-16'h0251,16'h0009,16'h0008,16'h0011,-16'h000d,16'h0010,16'h0013,-16'h002b,16'h000c,16'h001f,-16'h004a,16'h0021,16'h0018,16'h005c,-16'h0048,16'h0083,16'h0062,-16'h00a0,16'h0066,-16'h001a,16'h0008,-16'h0005,16'h0014,-16'h008e,16'h0050,16'h0004,16'h002f,16'h0019,-16'h004f,16'h002d,-16'h0007,-16'h0030,16'h003c,16'h0038,16'h0022,16'h0012,16'h005a,-16'h001f,16'h005a,-16'h000e,16'h0006,-16'h001d,16'h0021,-16'h0027,16'h0060,16'h005f,-16'h00a5,-16'h0025,16'h003b,-16'h002c,16'h0000,-16'h00a4,16'h0002,-16'h0007,16'h0071,16'h003a,16'h0004,16'h000e,-16'h0044,16'h0065,-16'h005c,-16'h0005,-16'h0019,16'h0058,-16'h01a0,16'h0000,-16'h0003,16'h0038,-16'h001c,16'h000e,16'h002e,-16'h0053,16'h0076,16'h0001,-16'h005f,16'h0021,16'h002f,16'h0043,-16'h0026,16'h003a,16'h006c,-16'h00b0,16'h0078,16'h0000,-16'h0017,16'h0044,16'h0013,-16'h017b,16'h0041,-16'h0012,16'h0030,16'h0000,-16'h0023,16'h001a,16'h0002,-16'h003e,16'h0049,16'h0046,16'h0045,-16'h0010,16'h0069,16'h0003,16'h003c,-16'h000c,16'h002d,16'h000e,16'h003b,16'h0013,16'h004d,16'h0069,-16'h00b8,-16'h0022,16'h0035,-16'h001c,16'h0000,-16'h00b2,-16'h0005,-16'h0011,16'h0032,16'h0030,16'h001a,-16'h000e,-16'h00b1,16'h0056,-16'h00a8,16'h000a,-16'h0009,16'h0036,-16'h00ac,-16'h0014,16'h0022,16'h0058,-16'h0009,-16'h0016,16'h0066,-16'h001c,16'h0087,16'h0007,-16'h00ac,16'h0002,16'h0038,16'h0023,16'h0008,-16'h0033,16'h0048,-16'h0046,16'h0057,16'h0011,16'h0028,16'h0061,16'h0000,-16'h01bf,16'h0065,-16'h0048,-16'h001a,-16'h0003,16'h001a,16'h0016,16'h0003,16'h0000,16'h0071,16'h002d,16'h0040,-16'h0027,16'h0062,16'h0014,16'h0044,16'h0005,16'h002b,16'h0010,16'h005c,16'h000b,16'h003d,16'h006c,-16'h00c9,-16'h0024,16'h000b,16'h0007,-16'h0007,-16'h00a2,16'h0012,16'h0012,16'h002d,16'h0016,16'h0022,-16'h000f,-16'h013b,16'h0069,-16'h0067,16'h0003,16'h0007,16'h003d,-16'h005e,-16'h0029,-16'h0011,16'h0037,16'h0001,16'h0004,16'h0077,-16'h002f,16'h0031,-16'h000d,-16'h00bb,-16'h001d,-16'h0012,16'h0031,16'h000f,-16'h005a,16'h002d,16'h0061,16'h005a,-16'h0007,16'h001c,16'h0066,16'h0001,-16'h0193,16'h005b,-16'h0040,-16'h0014,16'h000e,16'h001f,16'h0032,-16'h0013,-16'h002b,16'h0063,16'h0038,16'h003b,-16'h0022,16'h0083,-16'h0007,16'h002e,16'h0027,16'h002d,16'h0015,16'h004f,16'h0016,16'h0032,16'h0081,-16'h00a8,-16'h001d,16'h0038,16'h0020,16'h0028,-16'h00ba,16'h0000,16'h001e,-16'h002b,16'h0022,16'h003b,-16'h0026,-16'h0101,16'h0079,-16'h0007,-16'h0007,16'h0014,16'h002b,-16'h004b,16'h0002,16'h0001,16'h0023,-16'h0008,-16'h001a,16'h0096,-16'h003c,-16'h000d,-16'h001c,-16'h00a3,-16'h001f,-16'h004b,16'h0049,16'h001d,-16'h0060,16'h005c,16'h00bd,16'h004a,16'h000b,16'h0021,16'h0062,-16'h000c,-16'h013e,16'h0041,-16'h000d,-16'h001b,-16'h0002,16'h003b,16'h002e,-16'h004c,-16'h000f,16'h004a,-16'h000c,16'h0045,-16'h003a,16'h009a,-16'h0001,16'h0057,16'h0040,16'h0016,16'h000e,16'h0039,16'h0018,16'h002e,16'h005d,-16'h004e,-16'h0007,16'h0022,16'h001e,16'h000a,-16'h00cd,16'h000e,16'h002d,-16'h003d,16'h003b,16'h0014,-16'h0027,-16'h0088,16'h0061,16'h002c,16'h001a,16'h0003,16'h002c,-16'h0029,16'h0011,16'h0014,16'h002e,-16'h002d,-16'h003d,16'h0055,-16'h003d,-16'h0043,-16'h004e,-16'h0068,-16'h0029,-16'h00a5,16'h0034,-16'h000d,-16'h0043,16'h0066,16'h00dd,16'h003c,16'h0019,16'h002d,16'h006a,16'h0011,-16'h00cd,16'h002a,16'h000d,-16'h001c,16'h0001,16'h0036,16'h0060,-16'h0045,16'h000a,16'h0046,-16'h0074,16'h004f,-16'h0019,16'h0080,-16'h0009,16'h0068,16'h0050,-16'h0019,-16'h000f,16'h0003,16'h0028,16'h0000,16'h0048,-16'h0038,16'h0004,16'h001c,16'h0047,16'h0021,-16'h00b9,16'h0006,16'h001e,-16'h00b2,16'h004f,16'h0001,-16'h0018,16'h0012,16'h0054,16'h004a,16'h0036,-16'h0011,16'h001d,-16'h0023,-16'h0015,-16'h0020,16'h0002,-16'h002b,16'h0001,16'h0035,-16'h0026,-16'h0063,-16'h0039,-16'h0051,-16'h0032,-16'h0093,16'h002f,-16'h004b,16'h000f,16'h0094,16'h00b0,16'h0038,16'h0023,16'h003e,16'h0088,-16'h0006,-16'h0077,16'h0029,-16'h0020,16'h0014,16'h0011,16'h002a,16'h0054,-16'h0019,16'h0000,-16'h000c,-16'h00cd,16'h0077,-16'h0028,16'h005d,16'h0014,16'h000e,16'h0065,-16'h000b,-16'h002b,16'h0003,16'h000b,-16'h002c,16'h002a,-16'h0036,16'h0020,-16'h0008,16'h0053,16'h004a,-16'h0098,16'h000f,16'h0042,-16'h0103,16'h0057,16'h001e,-16'h0015,16'h008d,16'h0045,16'h006d,16'h0017,-16'h0006,16'h0029,-16'h002b,-16'h0040,-16'h0009,-16'h0028,-16'h0042,16'h000c,16'h0030,-16'h0031,-16'h007c,16'h0012,-16'h0026,16'h0013,-16'h0099,16'h002b,-16'h0044,16'h000f,16'h00a9,16'h004c,16'h0021,16'h001b,16'h0054,16'h008f,16'h0030,-16'h005c,16'h0028,-16'h000f,16'h0005,16'h0001,16'h001d,16'h0076,-16'h0012,-16'h0009,-16'h0036,-16'h00c2,16'h007a,-16'h001d,16'h0056,-16'h0008,-16'h0045,16'h006d,-16'h0025,-16'h0016,16'h000a,16'h001e,-16'h0022,16'h0002,-16'h0018,16'h000a,-16'h0018,16'h0067,16'h0039,-16'h0071,16'h000a,16'h001c,-16'h013b,16'h0049,16'h0007,-16'h0013,16'h0088,16'h005a,16'h007f,16'h0017,-16'h0011,16'h003b,-16'h0001,-16'h0030,-16'h002f,-16'h001f,-16'h002f,16'h003a,16'h0026,-16'h001a,-16'h0062,16'h0036,-16'h0020,16'h0009,-16'h0094,16'h0026,-16'h0020,16'h0000,16'h00d4,16'h001d,16'h003c,16'h001f,16'h0061,16'h008e,16'h0038,-16'h0044,16'h0040,16'h0022,16'h0017,16'h000a,16'h003f,16'h0070,-16'h0033,-16'h0011,-16'h0036,-16'h009b,16'h0043,16'h0010,16'h004b,-16'h000b,-16'h0082,16'h0086,16'h0022,-16'h0022,16'h000e,16'h003f,-16'h0056,-16'h0064,-16'h0026,-16'h0019,-16'h000d,16'h0026,16'h009e,-16'h006d,16'h005c,16'h0031,16'h000d,16'h0031,16'h0019,-16'h002c,16'h003d,16'h0051,-16'h005e,-16'h002a,-16'h0014,16'h0035,-16'h0057,16'h000a,16'h0085,16'h003c,-16'h0003,16'h006b,16'h002b,-16'h0028,16'h001c,16'h0035,-16'h0034,-16'h0015,16'h0026,-16'h000d,-16'h0002,16'h000e,16'h000a,16'h006d,16'h004d,16'h002e,-16'h004f,16'h0041,-16'h0002,16'h0049,-16'h003a,-16'h0035,16'h0058,-16'h001a,16'h000d,-16'h0061,-16'h0013,-16'h0043,-16'h0008,16'h0004,16'h0037,16'h0001,16'h0072,16'h0017,16'h0006,-16'h002b,16'h0029,16'h0002,16'h0006,16'h0034,-16'h0064,-16'h0036,-16'h0015,-16'h0004,16'h0013,16'h0012,16'h0074,-16'h0083,16'h0029,16'h003e,-16'h0011,16'h0030,-16'h0003,-16'h0016,16'h0036,16'h0040,-16'h0045,-16'h001b,-16'h001b,16'h0022,-16'h0020,-16'h0004,16'h008d,16'h0032,16'h0003,16'h007e,16'h002e,-16'h0039,16'h0001,16'h0035,-16'h003e,16'h0008,16'h001c,-16'h0010,-16'h0024,-16'h0018,-16'h0007,16'h0037,16'h0070,16'h002d,-16'h0062,16'h0038,-16'h001c,16'h005f,-16'h0067,-16'h0019,16'h0025,-16'h0015,16'h0069,-16'h001f,-16'h004f,-16'h0035,16'h0015,-16'h000a,16'h0044,16'h002d,16'h0049,16'h002b,16'h000b,16'h0000,16'h0022,-16'h000a,-16'h001b,16'h0035,-16'h0097,-16'h0010,-16'h0034,16'h0011,16'h001d,16'h001f,16'h003c,-16'h0097,16'h0008,16'h0077,-16'h0053,16'h0057,-16'h000c,16'h0033,-16'h000b,16'h002d,-16'h000e,-16'h000c,-16'h0038,16'h001f,-16'h0008,-16'h0032,16'h0050,16'h0018,-16'h000b,16'h0089,16'h0005,-16'h0019,-16'h003d,16'h002b,-16'h001e,-16'h000d,-16'h000a,-16'h0020,-16'h0044,-16'h002f,16'h0005,16'h000f,16'h0077,16'h0032,-16'h0059,16'h0004,16'h0019,16'h0050,-16'h0090,-16'h0013,16'h0033,-16'h0016,16'h0077,16'h000d,-16'h0043,-16'h0018,16'h000c,-16'h0003,16'h0037,16'h0058,16'h0022,16'h0019,16'h0014,-16'h000b,16'h0034,-16'h000c,-16'h004a,16'h0046,-16'h00c6,16'h0004,-16'h003d,-16'h0011,16'h0002,16'h003e,-16'h0006,-16'h0074,-16'h001b,16'h0052,-16'h0038,16'h003c,-16'h0017,16'h0057,-16'h0022,16'h0001,-16'h002d,-16'h0021,-16'h003a,16'h0006,-16'h0025,-16'h003e,16'h002f,16'h001b,-16'h001d,16'h0096,16'h0010,-16'h001d,-16'h0021,16'h0028,-16'h0003,16'h000a,16'h0000,-16'h0046,-16'h003e,-16'h0013,16'h0005,-16'h0024,16'h0088,16'h0044,-16'h004e,16'h000c,-16'h0008,16'h0051,-16'h008f,-16'h0019,16'h0041,-16'h001b,16'h0086,-16'h0002,-16'h0044,-16'h000f,16'h001f,-16'h0008,16'h0025,16'h0042,16'h000f,16'h0033,-16'h0013,16'h0000,16'h0051,-16'h0033,-16'h0044,16'h0060,-16'h008e,16'h001f,-16'h0077,16'h0007,16'h0011,16'h0039,16'h0022,-16'h0050,-16'h0013,16'h0059,-16'h002d,16'h0056,-16'h000e,16'h002d,-16'h0040,16'h001e,-16'h003c,-16'h000c,-16'h004e,16'h003e,-16'h001e,-16'h0016,-16'h0052,16'h002a,-16'h0005,16'h0059,16'h0020,16'h0010,16'h0017,16'h0007,16'h0029,-16'h0004,16'h000a,-16'h002d,-16'h001e,16'h000a,16'h0025,-16'h0014,16'h0093,16'h0048,-16'h001e,16'h0030,16'h0025,16'h0055,-16'h00af,16'h0002,16'h003b,-16'h0009,16'h00a5,16'h000c,-16'h003c,16'h0023,16'h0039,-16'h0001,16'h0027,16'h0052,16'h0010,16'h003f,-16'h0002,-16'h001d,16'h0062,-16'h0031,-16'h001d,16'h0041,-16'h004e,16'h0000,-16'h007e,16'h0001,16'h001c,16'h0056,16'h000d,-16'h0009,-16'h002d,16'h001b,-16'h0023,16'h004c,-16'h0035,-16'h0002,-16'h001f,16'h0020,-16'h0068,-16'h001e,-16'h004d,16'h0018,-16'h0028,-16'h0023,-16'h00b6,16'h0038,16'h002c,16'h007a,16'h0007,-16'h000b,16'h0010,16'h000a,16'h0052,16'h0004,-16'h0004,-16'h0045,16'h0019,-16'h0009,16'h002f,-16'h0004,16'h0088,16'h002e,-16'h000f,16'h003b,16'h0028,16'h0028,-16'h00bb,16'h0002,16'h002b,16'h0007,16'h0075,-16'h0031,-16'h0050,16'h0041,16'h0040,-16'h000a,-16'h0012,16'h0053,16'h0012,16'h003f,-16'h0012,16'h0000,16'h004e,-16'h0040,-16'h002e,16'h006a,-16'h0007,16'h000a,-16'h005a,-16'h0001,-16'h0001,16'h004a,16'h0000,16'h0043,-16'h0027,16'h000b,-16'h002e,16'h0059,-16'h001b,-16'h0056,-16'h0011,16'h0002,-16'h0066,-16'h0035,-16'h0014,16'h0019,-16'h0039,-16'h002c,-16'h0153,16'h003b,16'h0019,16'h007f,16'h0021,-16'h0023,-16'h0006,16'h0025,16'h005b,16'h0025,16'h001e,-16'h003c,-16'h0001,-16'h0019,16'h0040,16'h0010,16'h007e,16'h001b,16'h0028,16'h0044,16'h0000,16'h003f,-16'h0115,16'h002a,16'h000f,16'h000c,16'h001a,-16'h0023,-16'h0035,16'h0064,16'h0042,-16'h0013,16'h0004,16'h0038,16'h0024,16'h0046,-16'h000b,-16'h002f,16'h0037,-16'h0015,-16'h0009,16'h0037,16'h003a,-16'h0014,-16'h0064,-16'h0014,-16'h0016,16'h0026,-16'h000a,16'h0061,-16'h0027,-16'h0008,-16'h005c,16'h002a,-16'h004f,-16'h00a8,-16'h0018,-16'h0003,-16'h004e,-16'h003f,-16'h002e,16'h003a,-16'h0031,-16'h001c,-16'h0133,16'h004b,-16'h0012,16'h006f,16'h0009,-16'h0004,-16'h0018,16'h0022,16'h0055,16'h0011,16'h0008,-16'h0019,16'h002a,-16'h000e,16'h005b,-16'h0003,16'h0077,-16'h0006,16'h003b,16'h001e,-16'h001a,16'h003d,-16'h016c,16'h0006,16'h0009,16'h0057,-16'h0002,-16'h0019,-16'h002e,16'h0074,16'h002a,16'h0010,16'h0014,-16'h0036,16'h0031,16'h0021,-16'h000f,-16'h002f,16'h004e,-16'h0018,-16'h0013,16'h0033,16'h005f,-16'h0006,-16'h0061,-16'h0015,-16'h0043,16'h0003,-16'h0003,16'h00a6,-16'h0016,-16'h0006,-16'h0078,16'h0002,-16'h0024,-16'h0086,16'h0009,-16'h0008,-16'h003e,-16'h0033,-16'h002a,16'h003f,-16'h0029,-16'h006b,-16'h0039,16'h0023,-16'h0034,16'h006d,-16'h0003,16'h000a,16'h0004,16'h0027,16'h0077,16'h000d,-16'h0017,-16'h0018,16'h0058,-16'h0017,16'h006b,-16'h0026,16'h0064,16'h0008,16'h0020,16'h0048,16'h0011,16'h0018,-16'h0197,16'h0005,16'h0004,16'h0051,-16'h003b,16'h000a,-16'h003a,16'h0084,-16'h0001,16'h0029,-16'h0023,-16'h0054,16'h0035,16'h0024,-16'h0037,-16'h0035,16'h002d,-16'h0005,-16'h0033,16'h003d,16'h0042,-16'h002a,-16'h0067,-16'h0001,-16'h0054,-16'h0008,16'h0019,16'h00a4,-16'h0034,-16'h000b,-16'h005e,-16'h0007,-16'h003a,16'h0022,-16'h0020,16'h0002,-16'h004e,-16'h000c,-16'h001f,16'h005a,16'h0001,-16'h0090,16'h0015,16'h004e,-16'h0021,16'h006b,-16'h0003,-16'h0001,-16'h0020,16'h0013,16'h007c,-16'h0009,-16'h0014,16'h0006,16'h003e,-16'h0010,16'h00a3,-16'h0020,16'h0064,-16'h0029,16'h0017,16'h0060,16'h0014,16'h0013,-16'h0119,16'h0014,16'h0005,16'h0041,-16'h006d,-16'h0010,-16'h002e,16'h008f,16'h0004,16'h0029,-16'h0023,-16'h0080,16'h001f,16'h0008,-16'h0037,-16'h001e,16'h0025,-16'h0005,-16'h000a,16'h0037,16'h0026,-16'h0023,-16'h0069,-16'h0018,-16'h0058,16'h001e,16'h002c,16'h00a7,-16'h0023,-16'h0012,-16'h0045,16'h0000,-16'h002e,16'h004a,-16'h0038,16'h0026,-16'h0046,-16'h000f,16'h0000,16'h006f,16'h0028,-16'h0070,16'h0043,16'h0018,-16'h0024,16'h0055,-16'h0006,-16'h000b,-16'h002a,16'h0020,16'h007a,16'h0011,-16'h0021,-16'h0006,16'h0002,-16'h0004,16'h00c2,-16'h001a,16'h0066,16'h0007,16'h0013,16'h001c,-16'h0002,16'h0013,-16'h00c1,-16'h0010,16'h001e,16'h0027,-16'h00a4,-16'h000c,-16'h0028,16'h0097,16'h0000,16'h0026,16'h0008,-16'h0051,16'h004f,-16'h0004,-16'h0019,-16'h0039,16'h000c,16'h0000,16'h001f,-16'h001c,16'h0043,-16'h0009,-16'h0056,16'h000a,-16'h0035,16'h0026,16'h001e,16'h0081,-16'h0007,-16'h0019,-16'h0036,16'h000e,-16'h0047,16'h008f,-16'h0049,16'h002a,-16'h002b,-16'h0006,-16'h0001,16'h004a,16'h004e,-16'h0026,16'h0041,-16'h0001,-16'h0040,16'h0071,16'h0004,-16'h000c,-16'h0038,16'h0024,16'h0061,16'h0000,-16'h0030,-16'h0018,-16'h006b,16'h0018,16'h00eb,-16'h0029,16'h0086,16'h0004,16'h0017,16'h002b,16'h0000,16'h0033,-16'h0048,-16'h0021,16'h0012,16'h000e,-16'h008f,-16'h0025,16'h0010,16'h00a7,16'h0004,16'h0028,-16'h0008,-16'h0016,16'h0054,-16'h0005,16'h0006,-16'h0009,16'h0024,16'h000a,16'h0030,-16'h000f,16'h0032,16'h000f,-16'h008a,16'h0006,-16'h004d,16'h0003,16'h0021,16'h0072,-16'h0015,-16'h0007,-16'h0050,16'h0006,-16'h0032,16'h0061,-16'h0047,16'h0022,-16'h0044,16'h0000,16'h0020,16'h0057,16'h0072,16'h0030,16'h002e,-16'h000f,-16'h001c,16'h005f,-16'h000f,-16'h0011,16'h0004,-16'h0004,16'h0067,-16'h0021,-16'h0051,-16'h002e,-16'h008e,16'h0038,16'h00ed,16'h0005,16'h0083,16'h000a,16'h0012,16'h000c,16'h0010,16'h003e,-16'h0024,16'h000c,16'h001c,16'h0018,-16'h007d,-16'h000d,16'h0037,16'h007c,16'h0004,16'h0003,-16'h000d,16'h0033,16'h0057,-16'h0012,16'h0034,-16'h001a,16'h0000,-16'h001c,-16'h0006,-16'h0003,16'h0033,16'h0014,-16'h009d,16'h0000,-16'h002a,-16'h0002,16'h0026,16'h005e,-16'h0007,-16'h000d,-16'h0047,-16'h0022,-16'h0034,16'h002a,-16'h000f,16'h0050,-16'h003f,-16'h000e,16'h001e,16'h0030,16'h00ab,16'h0049,16'h003e,-16'h0008,16'h000c,16'h007d,16'h001b,-16'h002b,16'h0028,-16'h0027,16'h0063,-16'h0016,-16'h0039,-16'h001e,-16'h0089,16'h0019,16'h00c8,16'h0038,16'h009d,16'h000c,16'h0017,16'h000a,-16'h0003,16'h000a,-16'h0030,16'h0000,-16'h0004,16'h001a,-16'h0061,16'h000f,16'h0041,16'h0088,16'h0027,16'h0008,-16'h001c,16'h0066,16'h0077,-16'h000a,16'h0010,16'h0002,16'h0000,-16'h0007,16'h0011,16'h000b,16'h0027,16'h005f,-16'h009c,16'h0000,-16'h0030,16'h0006,16'h0024,16'h0028,16'h0010,-16'h000c,-16'h000b,-16'h003d,-16'h0040,-16'h0073,16'h003f,16'h0059,16'h0002,16'h0000,16'h0014,16'h002e,16'h0096,16'h0055,16'h004e,16'h001f,16'h001b,16'h0065,16'h0022,16'h0003,16'h0018,-16'h0018,16'h003a,-16'h001c,-16'h0023,-16'h0045,-16'h0034,-16'h0025,16'h00ca,16'h0024,16'h0097,16'h0041,16'h000b,16'h0015,16'h0006,16'h0002,-16'h0013,-16'h0006,-16'h001c,16'h0028,-16'h003a,16'h002e,16'h002c,16'h0078,16'h0014,16'h000c,-16'h005d,16'h0055,16'h008c,-16'h0034,-16'h0005,-16'h0014,16'h0000,-16'h001e,16'h001b,16'h0026,16'h002a,16'h006a,-16'h00a9,-16'h0001,16'h0001,16'h003c,16'h001a,16'h0001,16'h0018,-16'h0007,16'h0007,-16'h001b,-16'h001f,-16'h0099,16'h0046,16'h0086,16'h0015,-16'h0009,16'h0006,16'h0033,16'h006e,16'h0063,16'h0045,16'h000d,-16'h0008,16'h006b,16'h0013,-16'h001c,-16'h0045,-16'h0002,16'h0006,16'h000a,-16'h0017,-16'h0011,16'h0036,-16'h0095,16'h00a8,16'h0045,16'h0072,16'h0056,16'h001b,16'h000b,16'h0009,16'h0000,-16'h0018,-16'h000d,16'h0007,16'h0053,-16'h0042,16'h003a,16'h000f,16'h005a,16'h0000,16'h0023,-16'h0040,16'h0044,16'h008b,-16'h001c,16'h0012,-16'h002c,16'h0005,-16'h0007,16'h001e,16'h001f,16'h0007,16'h0059,-16'h00a1,16'h0019,-16'h000f,16'h003f,16'h0027,-16'h003d,-16'h0009,-16'h0011,16'h0071,-16'h0023,16'h000c,-16'h0068,16'h0049,16'h007d,16'h0010,16'h0003,-16'h001b,16'h001e,16'h001e,16'h004c,16'h004b,16'h000f,-16'h0037,16'h0068,16'h002b,-16'h0028,-16'h00a4,16'h0007,-16'h0030,16'h0018,-16'h0010,16'h0012,16'h001b,-16'h005d,16'h008a,16'h005d,16'h0093,16'h001a,16'h001d,-16'h0021,16'h001e,16'h004b,16'h0002,16'h0002,-16'h0001,16'h005c,-16'h004d,16'h003f,16'h0016,16'h0041,16'h0018,16'h0035,-16'h0049,16'h0000,16'h005a,-16'h000f,16'h0014,-16'h002c,-16'h0003,-16'h0011,-16'h0020,16'h0029,-16'h0009,16'h0061,-16'h0094,16'h0002,16'h0010,16'h001e,16'h0032,-16'h002e,-16'h000a,16'h0008,16'h0079,16'h001a,16'h0024,-16'h0013,16'h0075,16'h0099,16'h0009,16'h0028,-16'h0014,16'h002d,-16'h0086,16'h0054,16'h002a,16'h000a,-16'h003a,16'h0035,16'h0031,-16'h000e,-16'h0095,16'h0010,-16'h002d,16'h0015,-16'h001c,16'h0017,16'h0009,16'h000f,16'h008b,16'h0062,16'h0069,16'h0002,16'h002c,-16'h0022,16'h0032,16'h005a,16'h0029,16'h0001,-16'h0016,16'h0073,-16'h0037,16'h0063,16'h001d,16'h0054,16'h0013,16'h0020,-16'h0029,16'h0005,16'h0051,16'h000c,16'h0031,-16'h0021,16'h000b,-16'h0018,16'h0004,16'h001f,-16'h0021,16'h003c,-16'h0082,-16'h0007,16'h0010,-16'h0006,16'h0019,-16'h0040,16'h0003,-16'h000d,16'h0075,16'h001d,16'h0018,-16'h001b,16'h004a,16'h0087,-16'h001e,16'h0016,-16'h0005,16'h004f,-16'h017d,16'h0038,16'h001e,-16'h0012,-16'h0025,16'h0010,16'h002e,-16'h0013,-16'h005a,16'h0006,-16'h0040,16'h0004,-16'h002c,16'h0015,-16'h000d,16'h0059,16'h0093,16'h0000,16'h0067,-16'h0032,16'h000f,-16'h0029,16'h003f,16'h0033,16'h003b,-16'h0023,-16'h000f,16'h0034,-16'h0009,16'h0048,16'h000c,16'h003d,16'h0022,16'h000a,-16'h002f,-16'h0003,16'h005d,16'h000e,16'h0040,-16'h001a,16'h001b,-16'h001e,16'h000e,-16'h0002,-16'h0049,16'h0047,-16'h0074,-16'h001e,-16'h0009,-16'h0022,16'h0024,-16'h0047,16'h0000,-16'h0035,16'h005f,16'h000d,16'h002a,-16'h0005,16'h000e,16'h0078,-16'h0038,-16'h000f,-16'h000a,16'h003f,-16'h022d,16'h001d,-16'h0009,16'h000b,-16'h002f,16'h0017,16'h0009,-16'h0002,16'h0000,-16'h0002,-16'h007d,16'h0014,-16'h000c,16'h003b,-16'h003a,16'h0069,16'h0089,-16'h0086,16'h006c,-16'h0044,-16'h0007,-16'h0002,16'h0030,-16'h0036,16'h002c,16'h0008,-16'h0015,16'h0020,-16'h0016,16'h0026,16'h0019,16'h0029,16'h001e,16'h001e,16'h0028,-16'h0028,16'h0042,16'h0007,16'h0023,-16'h0011,16'h002e,-16'h000b,16'h004c,-16'h000f,-16'h0077,16'h0054,-16'h005b,-16'h0015,16'h0007,-16'h0006,16'h0021,-16'h0056,16'h000c,-16'h0017,16'h0058,16'h002e,16'h003d,-16'h0005,-16'h0013,16'h004d,-16'h004f,16'h0003,-16'h0003,16'h0044,-16'h01b4,-16'h001c,-16'h001f,16'h003b,-16'h0006,16'h001c,16'h002a,-16'h0016,16'h004e,-16'h0012,-16'h00c5,16'h0009,16'h001b,16'h0043,-16'h001e,16'h0038,16'h008b,-16'h009d,16'h006d,-16'h0034,16'h0000,16'h004c,16'h002b,-16'h0100,16'h0040,16'h0007,-16'h0004,16'h0020,-16'h001a,16'h0007,16'h001d,16'h0026,16'h0026,16'h003d,16'h0043,-16'h002c,16'h0066,-16'h0001,16'h0036,-16'h0012,16'h003a,-16'h000b,16'h0057,16'h0000,-16'h0093,16'h004e,-16'h0066,-16'h0019,-16'h0007,16'h002b,16'h0016,-16'h008a,-16'h000e,-16'h0013,16'h000d,-16'h0003,16'h002e,-16'h0009,-16'h00ae,16'h005f,-16'h00a9,-16'h000b,-16'h0014,16'h002e,-16'h00cb,-16'h002e,-16'h001d,16'h002d,16'h0001,16'h000f,16'h0063,-16'h0042,16'h0070,16'h000f,-16'h00e7,-16'h0047,16'h003b,16'h0043,16'h0008,-16'h001d,16'h0062,-16'h0051,16'h007e,-16'h0050,16'h0014,16'h0061,16'h0009,-16'h017c,16'h0053,16'h0002,-16'h0050,16'h003f,-16'h001d,16'h0016,16'h0005,16'h002f,16'h004c,16'h0032,16'h0053,-16'h0036,16'h0069,16'h0009,16'h0037,16'h0001,16'h0023,16'h000d,16'h0055,16'h0036,-16'h008b,16'h006b,-16'h0063,16'h0005,16'h000c,16'h001b,16'h003b,-16'h00a6,16'h000f,16'h0009,-16'h0001,16'h0004,16'h0029,-16'h0011,-16'h0145,16'h0051,-16'h009a,-16'h000e,-16'h0010,16'h0030,-16'h006d,-16'h001f,-16'h0021,16'h0025,16'h0006,-16'h0005,16'h0080,-16'h0042,16'h0040,-16'h001c,-16'h00b5,-16'h002d,16'h0001,16'h0028,16'h0000,-16'h0053,16'h006b,16'h001f,16'h0053,-16'h0034,16'h0037,16'h006a,-16'h0002,-16'h01b4,16'h005c,16'h0017,-16'h002f,16'h000f,16'h003d,-16'h0004,-16'h001f,16'h0008,16'h0043,16'h0017,16'h005e,-16'h0020,16'h0079,16'h0017,16'h005e,16'h0023,16'h0018,16'h0022,16'h006a,16'h003b,-16'h0078,16'h005d,-16'h007f,-16'h001c,-16'h000a,16'h0033,16'h0052,-16'h00a5,16'h0006,16'h001b,-16'h002d,16'h002b,16'h003a,-16'h0018,-16'h0111,16'h0049,-16'h0025,-16'h000b,-16'h001a,16'h003f,-16'h0033,-16'h001a,16'h0009,16'h0010,-16'h0013,-16'h0014,16'h0079,-16'h0049,-16'h000c,-16'h0021,-16'h00a4,-16'h004b,-16'h002c,16'h0031,16'h0023,-16'h007c,16'h0054,16'h00c1,16'h0036,-16'h0045,16'h0059,16'h0060,16'h0019,-16'h0195,16'h002f,16'h000f,-16'h0003,16'h0041,16'h0027,16'h002a,-16'h0039,16'h0014,16'h004a,-16'h002c,16'h0056,-16'h003e,16'h007b,-16'h0036,16'h004d,16'h0050,16'h0019,16'h0021,16'h0054,16'h003c,-16'h0074,16'h0042,-16'h0059,-16'h0003,-16'h0008,16'h002f,16'h0032,-16'h00ac,16'h0014,16'h0011,-16'h0049,16'h0039,-16'h0001,-16'h0011,-16'h00b7,16'h0052,-16'h0016,16'h0014,-16'h0017,16'h0032,-16'h003c,-16'h0013,16'h0009,16'h0009,-16'h0008,-16'h0019,16'h0041,-16'h0019,-16'h0055,-16'h0035,-16'h006a,-16'h003f,-16'h0084,16'h0024,16'h0013,-16'h003c,16'h007e,16'h00b5,16'h0019,-16'h0024,16'h0049,16'h006e,16'h0023,-16'h010c,16'h002c,-16'h0006,16'h0006,16'h003c,16'h0028,16'h0048,-16'h0034,16'h0006,16'h003d,-16'h009c,16'h0095,-16'h0040,16'h0084,-16'h0016,16'h0050,16'h006c,16'h0019,-16'h0003,16'h000a,16'h001d,-16'h0087,16'h0028,-16'h002c,-16'h0002,-16'h0012,16'h004c,16'h003e,-16'h008f,16'h0022,16'h0043,-16'h0079,16'h0059,-16'h000d,-16'h001e,16'h0013,16'h0049,16'h0026,16'h000d,-16'h0009,16'h0026,-16'h001a,-16'h0028,16'h0014,16'h001c,-16'h0014,-16'h002b,16'h0000,-16'h0036,-16'h0065,-16'h0051,-16'h003d,-16'h0016,-16'h00d0,16'h001b,-16'h003b,16'h001c,16'h0068,16'h00ca,16'h0023,-16'h001f,16'h0059,16'h0085,16'h001e,-16'h00b6,16'h001a,16'h0000,16'h002e,16'h0050,16'h0043,16'h0044,-16'h0019,16'h0010,16'h0015,-16'h00b7,16'h0068,-16'h0020,16'h006e,-16'h0012,-16'h002a,16'h0040,-16'h0029,-16'h0005,16'h0006,16'h0032,-16'h0075,16'h0001,-16'h0029,-16'h001e,-16'h0033,16'h004e,16'h0056,-16'h0093,16'h0012,16'h002f,-16'h00d5,16'h0053,-16'h001a,-16'h000d,16'h0091,16'h0035,16'h0061,-16'h0013,-16'h000d,16'h003e,-16'h002d,-16'h002c,-16'h000f,16'h000f,-16'h0023,16'h000e,16'h002c,-16'h003a,-16'h006d,-16'h000f,-16'h002e,-16'h000c,-16'h00b7,16'h0038,-16'h0030,16'h001d,16'h00aa,16'h0074,16'h0004,-16'h0034,16'h005d,16'h0091,16'h0023,-16'h008c,16'h0026,16'h0009,16'h002c,16'h004b,16'h0061,16'h0060,-16'h002f,-16'h0026,-16'h000a,-16'h00a1,16'h0075,-16'h0029,16'h0067,-16'h000c,-16'h0074,16'h004d,-16'h0028,-16'h0002,-16'h0010,16'h0035,-16'h0057,-16'h0026,-16'h001f,16'h0003,-16'h0035,16'h005f,16'h0068,-16'h0067,16'h001d,16'h0009,-16'h0138,16'h0050,-16'h000f,-16'h0016,16'h0099,16'h0034,16'h005d,16'h000c,-16'h0012,16'h0044,-16'h001f,-16'h0020,16'h0010,-16'h0026,-16'h001b,16'h0050,16'h0032,-16'h0036,-16'h006d,16'h000c,-16'h0029,16'h0009,-16'h0089,16'h0017,-16'h0028,16'h001e,16'h00d6,16'h0008,16'h0030,-16'h0026,16'h0066,16'h008b,16'h0026,-16'h004b,16'h002d,16'h000b,-16'h0003,16'h0069,16'h0021,16'h0065,-16'h004c,-16'h0039,-16'h0019,-16'h0075,16'h006c,16'h000c,16'h0069,-16'h0017,-16'h0092,16'h008c,-16'h0011,-16'h0024,16'h0008,16'h005a,-16'h0045,-16'h0064,-16'h002e,16'h0000,-16'h0012,16'h000f,16'h007b,-16'h0046,16'h0049,16'h0030,16'h0019,16'h002c,-16'h0024,-16'h0011,16'h0035,16'h0059,-16'h002d,-16'h002d,-16'h0023,-16'h0003,-16'h0017,16'h0004,16'h00a6,16'h002a,16'h0000,16'h008f,16'h0035,-16'h0038,16'h0004,16'h002d,-16'h002e,-16'h0008,-16'h0001,-16'h0028,16'h000d,-16'h0008,-16'h0014,16'h0052,16'h0046,16'h0048,-16'h002c,16'h0009,-16'h000b,16'h0048,-16'h003e,-16'h000f,16'h0030,16'h000d,16'h001c,-16'h0047,-16'h0001,-16'h0039,16'h0011,16'h0000,16'h0045,16'h0036,16'h004e,16'h001e,-16'h001f,-16'h000c,16'h003c,16'h0017,16'h001b,16'h0070,-16'h0064,-16'h0041,-16'h0029,16'h0018,16'h000b,16'h001e,16'h0041,-16'h0048,16'h0025,16'h004c,-16'h0023,16'h0025,-16'h0005,-16'h0001,-16'h000f,16'h0038,-16'h0026,-16'h0022,-16'h003d,-16'h000e,-16'h000f,-16'h0013,16'h0055,16'h0027,-16'h0019,16'h0094,16'h001d,-16'h0034,16'h0011,16'h0014,-16'h0039,-16'h0002,-16'h000a,-16'h0002,16'h0004,-16'h0029,-16'h0012,16'h000a,16'h0047,16'h0022,-16'h004a,-16'h0022,-16'h0012,16'h003a,-16'h0082,-16'h001c,16'h0024,16'h001c,16'h005e,16'h0012,-16'h0036,-16'h003a,16'h002c,16'h001b,16'h002a,16'h0030,16'h0023,16'h0025,-16'h0016,-16'h0012,16'h0040,16'h001c,-16'h002a,16'h0051,-16'h0092,-16'h001b,-16'h0057,16'h004a,16'h0002,16'h002c,16'h002b,-16'h0096,-16'h0002,16'h006c,-16'h0020,16'h0026,-16'h001e,16'h0056,-16'h0022,16'h0043,-16'h004a,-16'h002f,-16'h0033,16'h0015,-16'h000d,-16'h0046,16'h002f,16'h0017,-16'h002d,16'h007c,-16'h0007,-16'h0007,-16'h001c,16'h000f,-16'h001a,16'h0002,16'h0009,-16'h001b,-16'h0013,-16'h003f,-16'h001e,-16'h000e,16'h0038,16'h002c,-16'h006e,16'h000c,16'h0018,16'h003d,-16'h00a5,-16'h0022,16'h0026,-16'h000f,16'h0060,16'h003d,-16'h0049,-16'h003f,16'h001e,16'h0000,16'h0011,16'h0051,16'h0029,16'h0027,16'h0000,-16'h001f,16'h0049,-16'h0018,-16'h0033,16'h0025,-16'h0091,-16'h0017,-16'h006d,16'h0042,-16'h0017,16'h001d,16'h001e,-16'h0091,-16'h001e,16'h0051,-16'h000d,16'h0045,-16'h000b,16'h005b,-16'h0027,16'h0014,-16'h005f,-16'h0010,-16'h0024,-16'h000c,-16'h0010,-16'h0070,-16'h0002,16'h0004,-16'h001c,16'h0089,16'h001b,-16'h000d,16'h0000,16'h0018,-16'h0013,-16'h0001,-16'h002d,-16'h0006,-16'h0024,-16'h000b,-16'h0007,16'h0008,16'h006a,16'h0063,-16'h007a,16'h0008,-16'h0001,16'h0034,-16'h00c5,-16'h0022,16'h0020,16'h0024,16'h0086,16'h0028,-16'h005d,-16'h0025,16'h0011,16'h0005,16'h003e,16'h005e,16'h0021,16'h0035,-16'h0009,-16'h000d,16'h0058,-16'h001d,-16'h0039,16'h0024,-16'h003f,-16'h0018,-16'h0095,16'h004b,-16'h0019,16'h0037,16'h0024,-16'h0037,-16'h0013,16'h0038,-16'h001c,16'h0054,-16'h0028,16'h0019,-16'h003a,16'h0014,-16'h009c,-16'h001c,-16'h0036,16'h0015,-16'h001f,-16'h006b,-16'h0059,16'h002a,-16'h0010,16'h007a,16'h0006,-16'h0023,-16'h0003,16'h001d,16'h0013,-16'h0021,-16'h0025,16'h0002,-16'h0019,-16'h0027,16'h0009,-16'h0017,16'h0051,16'h0041,-16'h004b,16'h0000,-16'h0002,16'h0031,-16'h00bf,-16'h000f,16'h0027,16'h0050,16'h0084,16'h000d,-16'h0078,-16'h0027,16'h0008,-16'h0009,16'h003b,16'h0059,16'h0042,16'h0064,-16'h000d,-16'h0007,16'h0042,-16'h0023,-16'h004a,16'h0036,-16'h0016,-16'h0016,-16'h0098,16'h005e,-16'h0017,16'h0042,16'h0024,-16'h000c,-16'h0033,-16'h000a,16'h000a,16'h0035,-16'h0017,-16'h000e,-16'h0031,16'h0021,-16'h00b3,-16'h002a,-16'h003c,16'h0012,-16'h003c,-16'h0049,-16'h00c5,16'h004d,16'h001c,16'h00c8,16'h0020,-16'h002b,16'h0004,16'h000e,16'h0044,-16'h0001,-16'h0007,-16'h0031,16'h0017,-16'h001e,-16'h0010,16'h0011,16'h004f,16'h0028,16'h0008,16'h0010,16'h0012,16'h0042,-16'h00f2,-16'h0005,16'h001e,16'h0055,16'h0072,16'h001d,-16'h0058,-16'h0008,16'h0047,-16'h0012,16'h0033,16'h0027,16'h0034,16'h0055,-16'h0033,-16'h000a,16'h0038,-16'h0026,-16'h0050,16'h003b,16'h002e,-16'h0020,-16'h006b,16'h0043,16'h000d,16'h0039,16'h0002,16'h0054,-16'h0032,-16'h0008,-16'h0026,16'h003f,-16'h0013,-16'h00a9,-16'h0019,16'h0034,-16'h00c5,-16'h001c,-16'h005e,16'h002c,-16'h0020,-16'h0029,-16'h0119,16'h0040,16'h0006,16'h00a9,16'h0025,-16'h0020,-16'h0025,16'h0053,16'h003b,16'h000c,-16'h001e,-16'h0023,16'h001c,-16'h003a,16'h000a,16'h001e,16'h003f,16'h0002,16'h002f,16'h002a,16'h001f,16'h0052,-16'h014d,16'h0013,16'h003e,16'h0067,16'h0045,16'h0003,-16'h004c,16'h0034,16'h0055,-16'h001d,16'h0032,-16'h0024,16'h0031,16'h0025,-16'h001a,16'h0003,16'h0048,-16'h0023,-16'h003e,16'h0030,16'h004d,-16'h0030,-16'h0051,16'h003f,-16'h0006,16'h002f,16'h001d,16'h0081,-16'h0025,-16'h0014,-16'h005e,16'h0026,-16'h001e,-16'h00e0,-16'h0003,-16'h0004,-16'h008b,-16'h0042,-16'h0050,16'h003a,-16'h002e,-16'h004f,-16'h00a8,16'h002e,16'h0003,16'h00aa,16'h0034,-16'h000f,-16'h0009,16'h005b,16'h003f,16'h0004,16'h000e,-16'h002b,16'h0058,-16'h0026,16'h0009,16'h0017,16'h0036,-16'h0036,16'h0032,16'h0029,16'h0034,16'h0029,-16'h0169,16'h0002,16'h000e,16'h0096,16'h0005,16'h0009,-16'h0044,16'h006a,16'h003c,16'h0009,16'h003a,-16'h004e,16'h0020,16'h0016,-16'h0028,-16'h0007,16'h0034,-16'h0001,-16'h0034,16'h0006,16'h0050,-16'h0045,-16'h0027,16'h001f,-16'h0032,16'h0026,16'h0018,16'h0072,-16'h0028,-16'h002e,-16'h0084,16'h0009,-16'h0022,-16'h005c,-16'h0022,16'h0002,-16'h0086,-16'h0029,-16'h0046,16'h003d,16'h0005,-16'h0094,16'h0004,16'h0027,-16'h0017,16'h009a,-16'h001d,16'h0010,-16'h0007,16'h002a,16'h005f,16'h0004,-16'h000b,-16'h0003,16'h007d,-16'h0015,16'h0006,-16'h0006,16'h001d,-16'h0035,16'h0011,16'h001c,16'h000d,16'h0025,-16'h0138,-16'h0010,16'h0018,16'h0090,-16'h0038,16'h0018,-16'h003f,16'h009c,16'h0001,-16'h0005,16'h003a,-16'h005b,16'h0012,-16'h0010,-16'h0019,-16'h0001,16'h002e,-16'h0015,-16'h0009,16'h0018,16'h002c,-16'h0046,-16'h0013,16'h001c,-16'h0030,16'h000a,16'h0036,16'h0079,-16'h003b,-16'h0020,-16'h0083,16'h0009,-16'h0036,16'h003f,-16'h002b,16'h0027,-16'h0084,-16'h0016,-16'h0040,16'h0069,16'h0004,-16'h0075,16'h003c,-16'h0007,-16'h0043,16'h0074,16'h0000,-16'h0002,-16'h0029,16'h000a,16'h008b,16'h0013,16'h0001,-16'h000f,16'h0039,-16'h0017,16'h0040,-16'h0020,16'h001d,-16'h002e,16'h0022,16'h0040,16'h0008,16'h001e,-16'h00bf,-16'h001e,16'h0026,16'h0081,-16'h0084,16'h000a,-16'h0047,16'h00ba,-16'h0025,16'h000f,16'h0033,-16'h0051,16'h0021,-16'h001d,-16'h0035,-16'h0005,16'h0021,-16'h0010,16'h000b,16'h000d,16'h0034,-16'h0039,16'h0008,16'h0011,-16'h001d,16'h0025,16'h003c,16'h005e,-16'h002c,-16'h002d,-16'h0056,16'h000e,-16'h003e,16'h0096,-16'h002f,16'h0038,-16'h002a,-16'h0010,-16'h002d,16'h004d,16'h002d,-16'h003b,16'h0037,16'h000f,-16'h0039,16'h0065,16'h0007,-16'h000c,-16'h001f,16'h0015,16'h0081,-16'h000e,-16'h0009,-16'h0016,-16'h0025,-16'h0013,16'h0075,-16'h0014,16'h0029,-16'h0027,16'h002f,16'h002a,-16'h0013,16'h0045,-16'h0075,-16'h0013,16'h0017,16'h005f,-16'h00a4,16'h0003,-16'h0043,16'h00d5,-16'h000a,16'h0029,16'h001a,-16'h0010,16'h002f,-16'h0020,-16'h0008,-16'h000f,16'h003f,-16'h001a,16'h002f,16'h000b,16'h0036,-16'h0007,-16'h0008,16'h0019,-16'h0015,16'h001a,16'h0034,16'h0052,-16'h0034,-16'h0030,-16'h003c,16'h000a,-16'h004f,16'h0097,-16'h0048,16'h0034,-16'h0015,-16'h000d,-16'h000e,16'h0057,16'h0061,-16'h0033,16'h0045,16'h0000,-16'h0012,16'h007e,-16'h000a,16'h0003,-16'h001e,16'h000a,16'h0059,-16'h003f,-16'h0023,-16'h003e,-16'h008a,16'h0034,16'h00b9,-16'h0022,16'h0021,-16'h001c,16'h0021,16'h0021,-16'h0048,16'h0033,-16'h001d,-16'h000e,16'h0014,16'h0062,-16'h007d,-16'h0007,16'h0008,16'h00d4,16'h0013,16'h0033,16'h002d,16'h0000,16'h0030,-16'h0028,16'h000e,-16'h0006,16'h0016,-16'h000f,16'h0019,16'h0001,16'h0009,-16'h0001,16'h0002,16'h001e,-16'h000d,16'h0011,16'h0043,16'h0065,-16'h0015,-16'h000d,-16'h001a,-16'h0003,-16'h003f,16'h0067,-16'h0040,16'h005a,-16'h004b,-16'h000d,16'h0006,16'h0051,16'h0074,16'h0018,16'h0043,-16'h0015,16'h0000,16'h0088,-16'h000c,-16'h0023,16'h0013,-16'h0016,16'h006f,-16'h003a,-16'h0044,-16'h004a,-16'h0085,16'h0069,16'h00c5,16'h0013,16'h0027,16'h0015,16'h0003,-16'h0005,-16'h0043,-16'h000c,-16'h0016,-16'h0029,16'h0017,16'h0074,-16'h006d,16'h0010,16'h0036,16'h00e7,16'h0023,16'h002b,16'h000d,16'h0053,16'h0059,-16'h002c,16'h002f,-16'h001a,16'h0018,16'h0000,16'h0000,16'h000b,-16'h002a,16'h0039,-16'h0016,16'h0013,-16'h0007,16'h0003,16'h0029,16'h0061,16'h0005,-16'h0033,-16'h002f,-16'h001a,-16'h0040,-16'h0018,-16'h000c,16'h004d,-16'h0054,-16'h000a,-16'h000b,16'h0045,16'h0065,16'h0020,16'h0037,16'h0008,16'h0010,16'h008a,-16'h0019,-16'h0008,16'h0027,-16'h002c,16'h0034,-16'h0045,-16'h0023,-16'h0034,-16'h0051,16'h0046,16'h00ca,16'h0024,16'h0021,16'h0029,-16'h0021,-16'h001c,-16'h0038,-16'h002d,-16'h0027,-16'h0008,-16'h0007,16'h0053,-16'h0053,16'h0046,16'h0026,16'h00d5,-16'h0003,16'h0013,-16'h0008,16'h0061,16'h004b,-16'h002c,16'h0021,-16'h001d,16'h001b,-16'h0009,16'h0022,16'h0025,-16'h0075,16'h001e,-16'h0026,16'h000c,-16'h0012,16'h002a,16'h0045,16'h0028,16'h001d,-16'h0041,-16'h0018,-16'h0033,-16'h0041,-16'h00cc,16'h0020,16'h005b,-16'h001c,-16'h0002,16'h000a,16'h0038,16'h006e,16'h0042,16'h0067,16'h000c,16'h0038,16'h0090,16'h000c,16'h0008,16'h0015,-16'h0020,16'h0007,-16'h0037,-16'h002b,-16'h0016,-16'h000f,-16'h0030,16'h00bb,16'h001c,16'h0053,16'h003c,-16'h0007,16'h0007,-16'h000a,-16'h003a,-16'h0035,-16'h0030,-16'h001e,16'h006f,-16'h003f,16'h003c,16'h0027,16'h00d0,16'h000c,-16'h0013,-16'h0013,16'h0041,16'h005a,-16'h001c,16'h0035,-16'h0012,16'h0017,16'h0000,16'h003e,16'h0009,-16'h008f,16'h0036,-16'h0052,16'h000a,16'h0007,16'h004a,16'h0043,-16'h0009,16'h001e,-16'h003e,16'h0030,-16'h0014,-16'h0040,-16'h0098,16'h003c,16'h005e,16'h0012,-16'h0004,16'h000b,16'h0028,16'h0040,16'h0048,16'h0067,-16'h0001,-16'h0008,16'h0071,16'h0016,-16'h0019,-16'h002d,-16'h0009,-16'h003d,-16'h001a,-16'h0011,16'h0028,16'h0023,-16'h00b5,16'h00bc,16'h001d,16'h004a,16'h002b,16'h0028,-16'h0003,16'h0002,-16'h000a,16'h0003,-16'h0005,-16'h0037,16'h0066,-16'h001a,16'h004c,16'h000d,16'h009c,-16'h001b,-16'h0025,-16'h0026,16'h0042,16'h0055,-16'h0023,16'h0028,-16'h0018,16'h0001,-16'h0009,16'h0018,16'h002b,-16'h00b7,16'h005d,-16'h0043,16'h0001,-16'h0003,16'h005e,16'h004b,-16'h0036,16'h001a,-16'h003c,16'h0086,16'h0000,-16'h0003,-16'h004b,16'h0035,16'h0064,16'h0013,-16'h0003,-16'h0011,16'h0039,-16'h0009,16'h0047,16'h0050,16'h000e,-16'h0009,16'h0069,16'h001c,-16'h0015,-16'h007e,16'h0011,-16'h0051,16'h0026,-16'h0019,16'h000e,16'h003d,-16'h0073,16'h00be,16'h004a,16'h004a,16'h0004,16'h000e,-16'h001e,-16'h001c,16'h001e,16'h0000,16'h0001,-16'h003c,16'h009b,16'h0007,16'h0033,16'h0029,16'h0097,-16'h000c,-16'h0013,-16'h002c,16'h000f,16'h004e,-16'h0021,16'h001a,-16'h0020,-16'h0003,-16'h0024,-16'h0016,16'h0022,-16'h00d7,16'h0040,-16'h0025,-16'h0014,16'h0012,16'h004b,16'h0045,-16'h0031,16'h0021,-16'h0030,16'h007d,-16'h0003,-16'h001b,-16'h001f,16'h0029,16'h0058,-16'h0001,16'h0003,-16'h000d,16'h0024,-16'h0074,16'h0052,16'h000b,16'h0028,-16'h0013,16'h0026,16'h003b,-16'h0012,-16'h0096,16'h002f,-16'h0055,16'h002e,-16'h000b,16'h001c,16'h0001,16'h001f,16'h00b8,16'h0042,16'h003c,-16'h0021,16'h000d,-16'h002d,-16'h0002,16'h0047,16'h002f,16'h0005,-16'h0031,16'h006a,16'h0035,16'h0031,16'h0011,16'h008a,16'h0006,16'h0017,-16'h0036,-16'h0022,16'h0058,-16'h0002,16'h0022,-16'h0011,16'h0000,-16'h0027,-16'h0010,16'h0027,-16'h0108,16'h0024,-16'h000a,16'h0000,16'h000c,16'h000d,16'h0036,-16'h002d,16'h0029,-16'h001f,16'h006f,16'h0010,-16'h0012,-16'h000a,16'h0037,16'h006d,16'h0025,16'h0029,-16'h0006,16'h0032,-16'h0156,16'h003c,-16'h000a,16'h0016,-16'h0009,16'h002e,16'h0030,-16'h000c,-16'h007c,16'h0000,-16'h004c,16'h0027,-16'h0027,16'h000f,-16'h0003,16'h006b,16'h00c3,-16'h0015,16'h0017,-16'h003f,16'h000c,-16'h002c,16'h0004,16'h0056,16'h0016,16'h000c,-16'h002b,16'h005d,16'h002d,16'h0028,-16'h0005,16'h005d,-16'h0001,16'h0027,-16'h0020,-16'h006d,16'h0086,16'h001f,16'h0027,-16'h000d,16'h0010,-16'h0029,-16'h0009,-16'h0003,-16'h0110,16'h002c,16'h0000,16'h0015,-16'h001e,16'h0001,16'h004c,-16'h002b,16'h001d,-16'h0029,16'h004e,16'h0045,-16'h0009,16'h001e,-16'h000a,16'h004a,16'h0007,16'h0011,-16'h0020,16'h0021,-16'h01eb,16'h0020,-16'h0007,16'h0012,-16'h0008,16'h0033,16'h0034,-16'h0011,-16'h002e,-16'h0011,-16'h0083,16'h0026,-16'h001e,16'h0023,-16'h0017,16'h0057,16'h00c8,-16'h0086,16'h0011,-16'h005f,-16'h000b,-16'h002f,16'h0007,16'h000e,16'h0026,16'h0026,-16'h002b,16'h0050,16'h0023,16'h001b,16'h000d,16'h006f,-16'h000b,16'h0026,16'h0007,-16'h0053,16'h008a,16'h001b,16'h001b,-16'h0007,16'h000b,-16'h0038,16'h0003,-16'h000f,-16'h0140,16'h002c,16'h0009,16'h0003,16'h0001,-16'h000a,16'h0032,-16'h0025,16'h0004,-16'h0013,16'h0026,16'h0019,16'h0009,16'h0008,-16'h004c,16'h004f,-16'h004d,-16'h0009,-16'h001e,16'h0030,-16'h019a,-16'h0003,-16'h0026,16'h0003,-16'h001e,16'h004a,16'h0028,-16'h0008,16'h005d,16'h000a,-16'h00b9,-16'h0015,-16'h0017,16'h0061,-16'h0002,16'h004b,16'h008d,-16'h00b5,16'h0009,-16'h0069,-16'h0006,-16'h0016,16'h0003,-16'h0059,16'h0012,16'h002e,-16'h0039,16'h0058,-16'h002a,16'h0006,16'h002f,16'h0060,16'h0043,16'h0042,16'h0043,-16'h0032,16'h007f,16'h001b,16'h0021,16'h0002,16'h0036,-16'h002d,16'h0037,16'h0019,-16'h013c,16'h0035,16'h0013,16'h000f,-16'h000f,16'h0021,16'h005b,-16'h0038,-16'h0003,-16'h0008,16'h0015,16'h001a,16'h0025,16'h0002,-16'h00b1,16'h006c,-16'h0098,-16'h0028,-16'h0008,16'h0017,-16'h00de,-16'h0035,-16'h0032,-16'h0011,16'h000a,16'h004f,16'h002e,-16'h000a,16'h0086,-16'h0013,-16'h00e2,-16'h005e,16'h0028,16'h005d,16'h0002,-16'h0008,16'h0094,-16'h0040,16'h0000,-16'h0066,16'h0004,16'h003f,16'h0012,-16'h00be,16'h000b,16'h0052,-16'h0074,16'h0037,-16'h0022,-16'h0007,-16'h0005,16'h004a,16'h001a,16'h0037,16'h0054,-16'h002c,16'h0058,16'h0001,16'h0058,-16'h0004,16'h003b,-16'h0015,16'h005b,16'h0038,-16'h013d,16'h0045,16'h0009,16'h000c,-16'h0017,16'h003a,16'h0064,-16'h0064,16'h0016,16'h0017,-16'h0023,16'h0003,16'h0032,-16'h0017,-16'h016e,16'h0060,-16'h00a4,-16'h001e,-16'h0016,16'h0011,-16'h006e,-16'h0010,-16'h001a,-16'h000c,16'h0016,16'h0036,16'h005b,-16'h0006,16'h006d,-16'h001c,-16'h0092,-16'h0085,16'h0019,16'h0058,16'h0019,-16'h0049,16'h007a,16'h001b,16'h0019,-16'h0076,16'h002d,16'h006f,16'h0029,-16'h013f,-16'h0003,16'h003e,-16'h004b,16'h004f,16'h0002,16'h0000,-16'h0017,16'h0032,16'h0014,16'h0042,16'h0060,-16'h0021,16'h007d,-16'h0013,16'h0081,16'h001e,16'h000f,16'h0001,16'h0043,16'h0039,-16'h0113,16'h0057,-16'h0005,16'h0007,16'h0004,16'h003a,16'h0066,-16'h00d8,16'h0022,16'h0032,-16'h002d,16'h000f,16'h0032,-16'h0001,-16'h0150,16'h0035,-16'h0076,-16'h0026,-16'h003a,16'h0037,-16'h0062,-16'h0011,-16'h0017,16'h0016,-16'h0003,16'h000d,16'h0054,-16'h0027,16'h000c,-16'h000c,-16'h0077,-16'h0044,-16'h0013,16'h004b,16'h0007,-16'h005b,16'h0095,16'h00a7,16'h0015,-16'h0053,16'h0035,16'h0044,16'h002b,-16'h0196,-16'h000e,16'h0030,-16'h0022,16'h004a,16'h000b,16'h0016,-16'h003b,16'h0011,16'h0034,-16'h0024,16'h006d,-16'h0031,16'h0097,-16'h0039,16'h007b,16'h0025,16'h0006,16'h0005,16'h0034,16'h003a,-16'h0101,16'h002d,-16'h0013,16'h0013,-16'h001d,16'h0022,16'h006a,-16'h00d9,16'h0033,16'h0044,-16'h004b,16'h0023,-16'h0003,16'h0022,-16'h00d1,16'h0024,-16'h0022,-16'h0014,-16'h0025,16'h003b,-16'h0047,-16'h0002,-16'h0013,16'h0002,16'h0008,-16'h0004,16'h002f,-16'h0025,-16'h004f,-16'h0014,-16'h003e,-16'h0039,-16'h007b,16'h0025,-16'h0028,-16'h002c,16'h009b,16'h00cb,16'h001d,-16'h0076,16'h0055,16'h005f,16'h0032,-16'h015a,-16'h001b,-16'h0003,-16'h000f,16'h0051,16'h002e,16'h000f,-16'h0036,16'h0002,16'h0029,-16'h0072,16'h0086,-16'h0030,16'h009a,-16'h0025,16'h0022,16'h003e,-16'h0004,16'h000d,16'h002c,16'h0012,-16'h00d8,-16'h0017,-16'h002a,-16'h0003,-16'h0034,16'h003e,16'h0075,-16'h00bc,16'h0045,16'h0056,-16'h006d,16'h0053,-16'h0039,-16'h000c,-16'h000b,16'h0025,16'h0024,-16'h0020,-16'h002d,16'h0046,-16'h0026,-16'h001b,-16'h003c,16'h002e,-16'h002b,-16'h0002,16'h0009,-16'h000a,-16'h0055,-16'h0045,-16'h0023,-16'h001d,-16'h00d1,16'h0011,-16'h0027,16'h0018,16'h0090,16'h00d2,16'h001d,-16'h0053,16'h0046,16'h0088,16'h0037,-16'h00c6,-16'h0044,-16'h0013,16'h0018,16'h0051,16'h003c,16'h000e,-16'h000b,-16'h000a,16'h0001,-16'h0077,16'h0090,-16'h000e,16'h0074,-16'h0014,-16'h0054,16'h0015,16'h000b,16'h000f,16'h0007,16'h000b,-16'h00b2,-16'h0012,-16'h005f,-16'h0013,-16'h002b,16'h0049,16'h0063,-16'h0077,16'h002a,16'h004b,-16'h00b5,16'h0054,-16'h0005,16'h0001,16'h006a,16'h000c,16'h0064,16'h0005,-16'h0031,16'h0048,-16'h0038,16'h0001,-16'h001b,16'h0022,-16'h0016,16'h002b,16'h0018,-16'h0036,-16'h0053,-16'h0032,16'h0000,-16'h001f,-16'h00ca,-16'h0003,-16'h003a,16'h0032,16'h00a5,16'h008a,16'h001e,-16'h0065,16'h002c,16'h00a0,16'h0024,-16'h009d,-16'h0035,-16'h0027,16'h004a,16'h005b,16'h0047,16'h0038,-16'h0034,-16'h003e,-16'h001c,-16'h0062,16'h0073,-16'h0029,16'h0069,-16'h000f,-16'h0074,16'h0011,-16'h001a,-16'h0001,16'h0018,16'h0036,-16'h009c,-16'h0039,-16'h0055,-16'h0034,-16'h005b,16'h005d,16'h0071,-16'h0057,16'h0024,16'h0029,-16'h00f5,16'h0056,16'h002d,-16'h0018,16'h00b6,16'h0005,16'h006f,16'h0012,-16'h003f,16'h0069,-16'h0021,16'h0000,-16'h001b,16'h0005,-16'h004f,16'h003e,16'h0000,-16'h0022,-16'h005c,-16'h0001,-16'h000b,16'h0022,-16'h00ac,16'h0031,-16'h0035,16'h0037,16'h00d7,16'h003a,16'h001a,-16'h003f,16'h0054,16'h009b,16'h001d,-16'h006a,-16'h001a,-16'h000b,16'h0026,16'h0075,16'h001b,16'h0069,-16'h006d,-16'h005c,-16'h0024,-16'h005a,16'h006b,-16'h0006,16'h0067,-16'h001a,-16'h008d,16'h0084,-16'h0037,-16'h0009,-16'h0011,16'h0043,-16'h0049,-16'h002e,-16'h003d,16'h0002,-16'h0049,16'h0002,16'h0088,-16'h0041,16'h0024,16'h0014,16'h0021,16'h0040,-16'h001f,-16'h0003,16'h0013,16'h003a,-16'h0022,-16'h002f,-16'h000f,-16'h0009,16'h000a,16'h0024,16'h0070,16'h0049,-16'h002e,16'h0080,16'h003b,-16'h0036,16'h0004,16'h0013,-16'h0025,-16'h0013,-16'h0033,-16'h0032,16'h0017,-16'h000c,-16'h0037,16'h0039,16'h0032,16'h003a,-16'h0066,16'h0011,16'h000f,16'h0058,-16'h0046,-16'h0024,16'h001b,-16'h0009,16'h0028,16'h0005,16'h0001,-16'h0057,16'h0018,-16'h0004,16'h0033,16'h005e,16'h0035,16'h002b,-16'h000d,-16'h0025,16'h0015,16'h002b,16'h0017,16'h006f,-16'h007d,-16'h0040,-16'h0025,16'h0033,-16'h0039,16'h0014,16'h0043,-16'h0063,16'h0016,16'h004a,16'h0000,16'h002c,-16'h0008,16'h0025,16'h0004,16'h003a,-16'h000c,-16'h0032,-16'h002e,-16'h0018,16'h000f,-16'h0023,16'h0000,16'h001e,-16'h0022,16'h0084,16'h0014,-16'h0022,-16'h000e,16'h0009,-16'h004c,-16'h0003,-16'h0040,-16'h0001,-16'h0017,-16'h0036,-16'h0036,16'h0003,-16'h0001,16'h0023,-16'h0078,16'h0001,16'h003a,16'h004e,-16'h0063,-16'h000d,16'h001a,16'h000a,16'h0045,16'h0043,-16'h0040,-16'h0044,16'h0037,-16'h0006,16'h0019,16'h003d,16'h0029,16'h001d,-16'h0005,-16'h0030,16'h0032,16'h001d,-16'h0001,16'h003d,-16'h0084,-16'h0012,-16'h0040,16'h0045,-16'h0018,16'h000a,16'h0021,-16'h007c,-16'h0014,16'h0033,-16'h0032,16'h003c,-16'h0018,16'h0055,-16'h0019,16'h0044,-16'h0046,-16'h0022,-16'h0015,16'h0006,-16'h0001,-16'h0092,-16'h0007,16'h0004,-16'h0020,16'h0082,16'h0007,-16'h0016,16'h0000,16'h0004,-16'h0036,16'h0002,-16'h001f,16'h001f,16'h0000,-16'h0025,-16'h001f,16'h001b,16'h001b,16'h004f,-16'h007f,16'h0004,16'h001e,16'h0055,-16'h0081,-16'h002c,16'h0020,16'h004e,16'h0047,16'h0048,-16'h0036,-16'h002a,16'h0018,16'h0011,16'h0023,16'h005c,16'h0002,16'h0030,16'h0023,-16'h001c,16'h0010,-16'h000c,-16'h0048,16'h0045,-16'h0041,-16'h003e,-16'h0052,16'h0046,-16'h0039,16'h001c,16'h002d,-16'h0073,16'h0010,16'h002c,-16'h0023,16'h001d,16'h0007,16'h004c,-16'h0045,16'h0037,-16'h0071,-16'h0026,-16'h0040,16'h001d,16'h0011,-16'h00a9,-16'h001e,-16'h000e,16'h0009,16'h005d,-16'h001b,-16'h0020,-16'h0005,16'h000e,-16'h001e,16'h0002,-16'h002f,-16'h000d,-16'h0019,16'h0000,-16'h000d,-16'h0010,16'h0040,16'h0041,-16'h005f,16'h0010,16'h0033,16'h002d,-16'h0092,-16'h002c,16'h0021,16'h005d,16'h0063,16'h0045,-16'h0065,-16'h0036,-16'h0003,16'h0009,16'h0034,16'h0061,16'h002e,16'h005a,16'h001a,-16'h002d,16'h0015,-16'h000c,-16'h004e,16'h003a,-16'h0035,-16'h001b,-16'h0077,16'h0054,-16'h002e,16'h0012,16'h001b,-16'h000f,16'h000c,16'h000c,-16'h0034,16'h0017,16'h0003,16'h001a,-16'h0031,16'h0035,-16'h00a1,-16'h0021,-16'h002d,16'h001a,-16'h0010,-16'h006f,-16'h008f,16'h0009,16'h0010,16'h0068,16'h0028,-16'h0018,16'h0011,16'h000e,16'h0025,-16'h0003,-16'h0028,16'h000d,-16'h001d,-16'h0019,16'h0015,16'h0001,16'h003a,16'h003d,-16'h003a,-16'h0009,16'h0018,16'h0042,-16'h00b5,-16'h0011,16'h001b,16'h0056,16'h0051,16'h0032,-16'h0074,-16'h0033,16'h0021,16'h0000,16'h0047,16'h0072,16'h0056,16'h0060,-16'h0010,-16'h0004,-16'h0007,-16'h000f,-16'h003a,16'h003f,16'h002a,-16'h0029,-16'h004d,16'h0056,-16'h0008,16'h0006,16'h0022,16'h002b,-16'h0013,-16'h000e,-16'h0006,16'h0033,16'h0006,-16'h002e,-16'h0029,16'h0035,-16'h008b,-16'h0018,-16'h004f,16'h0021,-16'h0032,-16'h004c,-16'h00ef,16'h0000,16'h0021,16'h0099,16'h0020,-16'h0034,16'h000b,16'h000d,16'h001f,-16'h0017,-16'h0035,-16'h0021,-16'h0019,-16'h002b,16'h0006,16'h000d,16'h001b,16'h0048,16'h0014,-16'h0008,16'h000b,16'h0042,-16'h00e8,-16'h0001,16'h0029,16'h007b,16'h0070,16'h0038,-16'h0061,-16'h0055,16'h003f,-16'h0011,16'h0044,16'h0039,16'h001f,16'h003d,16'h0006,-16'h0005,16'h0010,-16'h000d,-16'h004b,16'h002f,16'h0036,-16'h0033,-16'h0059,16'h006d,16'h0011,16'h0028,16'h000a,16'h007b,-16'h0042,-16'h0030,-16'h0019,16'h0010,-16'h0010,-16'h00b4,-16'h0026,16'h0026,-16'h006b,-16'h0017,-16'h0043,16'h000a,-16'h000d,-16'h0036,-16'h00d4,16'h0022,-16'h0006,16'h00b0,16'h0006,-16'h003b,-16'h000e,16'h002f,16'h0038,-16'h0029,-16'h000a,-16'h0035,16'h0038,-16'h001a,-16'h0028,16'h002d,16'h0017,-16'h002f,16'h002e,-16'h0002,16'h0011,16'h004c,-16'h010b,16'h0006,16'h0016,16'h0093,16'h003d,16'h0043,-16'h0043,-16'h004d,16'h0036,-16'h0012,16'h003c,-16'h0023,-16'h0006,16'h000e,-16'h0017,16'h000a,16'h0016,-16'h0002,-16'h0032,16'h0022,16'h004d,-16'h0052,-16'h0039,16'h0076,16'h002d,16'h0008,16'h0017,16'h006c,-16'h0020,-16'h002c,-16'h003a,16'h0015,-16'h0002,-16'h00b5,-16'h0024,16'h0024,-16'h006e,-16'h0016,-16'h003f,16'h001c,-16'h0007,-16'h0068,-16'h001a,16'h0034,16'h0007,16'h00a5,16'h000d,-16'h002b,-16'h0021,16'h003b,16'h004d,-16'h0026,-16'h0007,-16'h002d,16'h008f,-16'h005e,-16'h0029,16'h000b,-16'h000c,-16'h003b,-16'h0003,16'h0019,16'h001c,16'h004a,-16'h00ef,16'h0003,16'h0008,16'h00ab,16'h0002,16'h004a,-16'h004c,-16'h0023,16'h001f,-16'h002a,16'h005d,-16'h0056,16'h0017,-16'h000b,-16'h0019,-16'h0003,16'h0041,-16'h0032,-16'h0031,16'h0000,16'h0032,-16'h0065,-16'h0001,16'h0078,16'h0032,16'h0000,16'h0041,16'h005f,-16'h002e,-16'h0034,-16'h0027,16'h0002,16'h0007,-16'h0004,-16'h002a,16'h0017,-16'h0041,-16'h001b,-16'h0061,16'h0037,-16'h001b,-16'h008f,16'h0031,16'h003c,-16'h0016,16'h00a1,-16'h0019,-16'h001b,-16'h0029,16'h001b,16'h004b,-16'h001d,-16'h001f,-16'h000f,16'h0059,-16'h003b,-16'h003e,16'h0003,-16'h001f,-16'h0047,16'h0008,16'h0019,-16'h0003,16'h0023,-16'h0091,16'h0003,16'h000d,16'h00a1,-16'h004c,16'h0041,-16'h0069,-16'h001c,16'h000b,-16'h000a,16'h003d,-16'h0057,16'h0013,-16'h0014,-16'h0022,-16'h0006,16'h0051,-16'h0026,-16'h000e,16'h0002,16'h0015,-16'h003b,16'h0012,16'h004c,16'h0061,16'h0003,16'h002b,16'h0037,-16'h0022,-16'h002e,-16'h0022,16'h000b,-16'h000e,16'h0069,-16'h0032,16'h0032,-16'h0038,-16'h001d,-16'h0056,16'h003e,-16'h0017,-16'h005c,16'h003d,16'h0029,-16'h0022,16'h0078,-16'h002a,-16'h002c,-16'h0024,16'h0010,16'h0086,16'h0000,-16'h000d,16'h001d,-16'h0011,-16'h0021,-16'h0015,-16'h0004,-16'h002b,-16'h0019,16'h000b,16'h0032,16'h0000,16'h0008,-16'h0064,16'h0004,16'h0034,16'h0094,-16'h0096,16'h0024,-16'h0058,16'h0038,16'h0000,16'h001d,16'h0028,-16'h0056,-16'h0013,-16'h0038,16'h0001,16'h0005,16'h0060,-16'h0034,16'h0008,-16'h002d,16'h001c,-16'h002c,16'h0032,16'h0038,16'h0063,-16'h0002,16'h002a,16'h0030,-16'h001e,-16'h0038,-16'h002a,-16'h0009,-16'h0018,16'h009b,-16'h0045,16'h0042,-16'h0016,-16'h0018,-16'h0032,16'h0037,16'h000b,-16'h0041,16'h0045,16'h001f,-16'h0028,16'h0063,-16'h000f,-16'h001a,-16'h0033,-16'h001a,16'h0060,-16'h0050,16'h0000,-16'h0017,-16'h0065,16'h0029,-16'h0017,-16'h000c,-16'h004e,-16'h0029,16'h0026,16'h005a,-16'h000a,16'h0038,-16'h002e,16'h0006,16'h003d,16'h007d,-16'h0086,16'h000f,-16'h002d,16'h0026,16'h000d,16'h0008,16'h0049,-16'h001d,16'h0004,-16'h001b,16'h0009,16'h0025,16'h003c,-16'h001d,16'h0031,-16'h0025,16'h000c,-16'h003d,16'h005a,16'h0041,16'h0058,16'h000c,16'h0008,16'h003a,16'h000c,-16'h0047,-16'h001c,-16'h0017,-16'h0040,16'h0081,-16'h005a,16'h005f,16'h0001,16'h0006,-16'h0008,16'h0047,16'h002f,-16'h0039,16'h0056,16'h000f,-16'h0007,16'h0090,-16'h0010,-16'h0010,-16'h002a,16'h0014,16'h006b,-16'h0061,-16'h0017,-16'h002a,-16'h00a2,16'h0040,16'h0016,16'h0006,-16'h0054,-16'h002c,16'h0011,16'h0039,-16'h0001,16'h0000,-16'h0017,-16'h0011,16'h0041,16'h0085,-16'h005f,16'h000c,16'h0012,16'h0046,16'h0037,16'h001a,16'h003c,16'h0025,-16'h0004,-16'h0017,16'h0041,-16'h000e,16'h0038,-16'h0027,16'h001f,-16'h0002,-16'h002e,16'h0000,16'h0082,16'h0034,16'h006e,16'h0000,16'h001f,16'h0066,16'h000b,-16'h0013,-16'h0022,-16'h0038,-16'h0060,16'h0057,-16'h0045,16'h0061,-16'h0058,-16'h0008,-16'h000b,16'h0046,16'h004c,-16'h000f,16'h0047,16'h0009,16'h0025,16'h0089,-16'h0008,-16'h0013,16'h0036,-16'h0006,16'h0068,-16'h0055,-16'h000a,-16'h0023,-16'h008a,16'h0093,16'h0036,16'h000b,-16'h0061,-16'h0011,-16'h000f,16'h0007,-16'h003a,16'h0001,-16'h0012,-16'h0036,16'h0025,16'h0085,-16'h0036,16'h001b,16'h003c,16'h0051,16'h005a,16'h0011,16'h001e,16'h005c,16'h0010,-16'h002d,16'h002b,-16'h000c,16'h003c,-16'h0016,16'h0002,16'h0000,-16'h0059,16'h001e,16'h0096,16'h0031,16'h0056,16'h001f,16'h0027,16'h0027,16'h000e,-16'h001d,-16'h0037,-16'h0024,-16'h004e,-16'h0060,-16'h0018,16'h0060,-16'h0068,-16'h0004,-16'h0022,16'h002b,16'h0041,16'h0019,16'h0048,16'h0008,16'h0035,16'h007e,16'h0015,-16'h0018,16'h0035,-16'h0025,16'h002e,-16'h0058,-16'h002e,-16'h0023,-16'h0043,16'h005d,16'h0044,16'h0011,-16'h0074,-16'h000f,-16'h0041,-16'h0041,-16'h003f,-16'h003b,16'h0003,-16'h003e,16'h001b,16'h007d,-16'h003e,16'h0031,16'h0022,16'h0083,16'h0036,-16'h000d,16'h0013,16'h0040,16'h0034,-16'h0033,16'h0038,-16'h0020,16'h0021,-16'h001e,16'h002f,-16'h0002,-16'h0049,16'h0002,16'h0061,16'h0035,16'h006d,16'h0026,16'h002f,-16'h0012,16'h0019,-16'h0011,-16'h0015,-16'h002b,-16'h0072,-16'h00b1,16'h0000,16'h0044,-16'h0016,16'h000e,-16'h0037,16'h001c,16'h0046,16'h0029,16'h0041,-16'h0011,16'h0044,16'h0093,16'h0021,-16'h0019,16'h005d,-16'h000b,-16'h0020,-16'h002b,-16'h002d,-16'h002c,-16'h0019,-16'h004d,16'h0079,16'h002b,-16'h0072,-16'h0019,-16'h001f,-16'h0016,-16'h0023,-16'h0029,-16'h0029,-16'h0048,16'h000d,16'h007d,-16'h002c,16'h0031,16'h0036,16'h0089,16'h0010,-16'h001f,-16'h0019,16'h0039,16'h0049,-16'h0046,16'h002e,-16'h0024,16'h0028,-16'h0010,16'h0005,16'h0007,-16'h0068,16'h002e,16'h0066,16'h0024,16'h0039,16'h002d,16'h0025,-16'h0024,16'h0027,-16'h0024,16'h000c,-16'h000a,-16'h005a,-16'h005c,-16'h0004,16'h0030,16'h000c,16'h0009,-16'h0035,16'h0036,16'h0057,16'h0035,16'h0053,-16'h0008,16'h000b,16'h0075,16'h0034,-16'h000d,-16'h0014,16'h0010,-16'h0030,16'h0012,-16'h001c,-16'h0023,16'h0027,-16'h00d4,16'h0085,16'h002d,-16'h0080,-16'h0014,16'h0006,-16'h000f,-16'h0059,-16'h0032,-16'h0049,-16'h003f,-16'h000b,16'h007c,16'h002b,16'h0026,16'h0039,16'h0083,16'h001b,16'h0003,-16'h003e,16'h0018,16'h0058,-16'h0017,16'h0004,-16'h0018,16'h000e,-16'h0015,-16'h0005,16'h0034,-16'h0073,16'h001d,16'h004d,16'h0048,16'h0016,16'h003b,16'h0050,-16'h0031,16'h0024,-16'h000b,16'h003a,-16'h000e,-16'h006e,-16'h000b,16'h0038,16'h004c,16'h002d,-16'h0004,-16'h003c,16'h0006,16'h0018,16'h004b,16'h001b,16'h0027,-16'h0004,16'h004b,16'h0031,-16'h0027,-16'h0063,16'h0038,-16'h005b,16'h0032,-16'h000f,-16'h000a,16'h0009,-16'h0073,16'h0075,16'h005e,-16'h007f,-16'h003f,16'h0026,-16'h0014,-16'h0065,16'h000e,-16'h000b,-16'h0013,-16'h001b,16'h0083,16'h0039,16'h0031,16'h0043,16'h005d,16'h0013,16'h0008,-16'h0055,-16'h0031,16'h0075,-16'h000f,16'h000e,-16'h0014,16'h0028,-16'h0026,-16'h0044,16'h0017,-16'h008c,16'h0025,16'h0059,16'h0019,16'h0033,16'h005b,16'h0058,-16'h0046,16'h0039,16'h0000,16'h006a,16'h000f,-16'h006a,-16'h0016,16'h0051,16'h0046,16'h0020,-16'h0003,-16'h0038,16'h003b,-16'h0025,16'h003d,16'h000b,16'h003c,-16'h0008,16'h0051,16'h0048,-16'h001a,-16'h009c,16'h002b,-16'h0054,16'h0056,-16'h0021,-16'h000c,-16'h002a,16'h0048,16'h0088,16'h0050,-16'h0076,-16'h0030,16'h002d,-16'h003c,-16'h005e,16'h0025,16'h0012,-16'h000c,-16'h0022,16'h006d,16'h0050,16'h003c,16'h001d,16'h0056,16'h000b,16'h0023,-16'h0054,-16'h0059,16'h006a,-16'h0017,16'h0006,16'h0002,16'h002c,-16'h0036,-16'h0046,16'h002a,-16'h00d4,16'h0020,16'h006d,16'h001f,16'h0011,16'h0017,16'h005f,-16'h0041,16'h003e,-16'h0025,16'h0079,16'h0005,-16'h005c,16'h0004,16'h0057,16'h0051,16'h0028,16'h001b,-16'h0031,16'h0018,-16'h00ed,16'h0036,-16'h000c,16'h0033,16'h0005,16'h003d,16'h0032,-16'h0033,-16'h008a,16'h0017,-16'h0079,16'h002e,-16'h0039,16'h0011,-16'h0014,16'h0067,16'h0090,-16'h0024,-16'h0097,-16'h0035,16'h001c,-16'h001a,-16'h0029,16'h0022,-16'h0002,-16'h0004,-16'h003b,16'h003f,16'h004a,16'h001f,16'h0027,16'h006a,16'h0018,16'h001c,-16'h0010,-16'h0083,16'h0075,16'h000a,16'h0002,-16'h001e,16'h001e,-16'h003c,-16'h003f,16'h002d,-16'h010e,16'h0025,16'h0065,16'h0037,-16'h0013,16'h0013,16'h0060,-16'h0034,16'h0054,-16'h0007,16'h005e,16'h0005,-16'h0024,16'h000d,16'h001b,16'h0037,-16'h0002,16'h000a,-16'h002d,16'h0011,-16'h01d5,16'h000f,-16'h0019,16'h0001,16'h001f,16'h0036,16'h0037,-16'h0010,-16'h0053,16'h000d,-16'h0088,16'h0011,-16'h0025,16'h004e,-16'h0014,16'h0056,16'h008c,-16'h00b8,-16'h0097,-16'h004e,-16'h0003,-16'h0026,-16'h0025,16'h0014,-16'h000d,16'h0019,-16'h002d,16'h0059,16'h0039,16'h000f,16'h000f,16'h0058,16'h0000,16'h002a,-16'h000d,-16'h0066,16'h00a5,16'h0014,16'h0027,-16'h0009,16'h0018,-16'h004a,-16'h0023,16'h000a,-16'h014d,16'h0018,16'h003e,16'h0024,-16'h0012,16'h0014,16'h004e,16'h0000,16'h0026,-16'h000c,16'h002b,16'h001b,-16'h0020,-16'h0008,-16'h004c,16'h003c,-16'h001b,16'h000d,-16'h0035,16'h0033,-16'h019f,-16'h0002,-16'h0020,-16'h0021,16'h0001,16'h0069,16'h000a,-16'h0021,16'h004f,16'h000a,-16'h00a8,-16'h0024,-16'h000d,16'h0063,-16'h0010,16'h0057,16'h00a8,-16'h00aa,-16'h0090,-16'h007e,16'h0009,16'h0023,-16'h000e,-16'h000f,-16'h002d,16'h0037,-16'h004b,16'h006d,16'h0029,16'h0006,16'h001c,16'h004c,16'h0013,16'h0037,16'h001a,-16'h0029,16'h00ab,16'h0002,16'h003c,16'h0015,16'h001b,-16'h0031,16'h0006,16'h0018,-16'h0195,16'h0009,16'h001f,16'h003f,-16'h0003,16'h0012,16'h0070,-16'h000f,16'h0026,16'h000a,16'h0013,16'h0015,16'h001c,-16'h0008,-16'h00c1,16'h0036,-16'h007f,-16'h0024,-16'h0024,16'h000c,-16'h0109,16'h0000,-16'h0015,-16'h0014,16'h0013,16'h0095,16'h001b,-16'h000c,16'h0076,-16'h000a,-16'h007c,-16'h0067,16'h0023,16'h007f,16'h0008,-16'h0013,16'h008f,-16'h0078,-16'h0071,-16'h0064,16'h0010,16'h001d,-16'h001c,-16'h0044,-16'h002b,16'h005c,-16'h0064,16'h0039,-16'h0001,16'h0008,-16'h0009,16'h004d,16'h0032,16'h002f,16'h0034,16'h0006,16'h0080,16'h0006,16'h003f,16'h0017,16'h0039,-16'h0053,16'h0051,16'h0029,-16'h0182,16'h0033,16'h0023,16'h002f,-16'h000d,16'h001f,16'h0058,-16'h002f,16'h0033,16'h0010,-16'h000b,16'h0023,16'h000b,16'h0003,-16'h0193,16'h001c,-16'h00aa,-16'h001f,-16'h002d,-16'h000d,-16'h009a,-16'h003b,-16'h000e,-16'h0001,16'h001c,16'h0061,16'h000f,-16'h0027,16'h006f,-16'h003f,-16'h0026,-16'h004f,16'h0016,16'h0063,-16'h0001,-16'h0070,16'h00ac,16'h000b,-16'h0049,-16'h0057,16'h0034,16'h003d,16'h001b,-16'h00bb,-16'h0035,16'h0026,-16'h0053,16'h0038,-16'h0008,-16'h0001,-16'h003b,16'h003f,16'h0017,-16'h002c,16'h002b,-16'h0007,16'h0050,-16'h000b,16'h0063,16'h001d,16'h000a,-16'h0048,16'h0055,16'h003c,-16'h0143,16'h000c,16'h000d,16'h001e,-16'h001f,16'h004c,16'h0078,-16'h0084,16'h003a,16'h0044,-16'h0021,16'h0011,16'h0011,16'h0015,-16'h0163,16'h0003,-16'h0063,-16'h0035,-16'h001c,-16'h0007,-16'h0069,-16'h000f,16'h0006,-16'h000e,16'h000f,16'h002d,16'h001e,-16'h002a,16'h0018,-16'h0028,-16'h0018,-16'h005d,16'h0004,16'h0043,16'h0026,-16'h0096,16'h00a3,16'h006e,-16'h001c,-16'h0056,16'h002a,16'h004e,16'h0035,-16'h0124,-16'h004c,16'h0018,-16'h0033,16'h0036,16'h0008,-16'h0023,-16'h005c,16'h0017,16'h0001,-16'h0036,16'h005a,16'h000b,16'h0072,-16'h002a,16'h0064,16'h0031,-16'h0021,-16'h0045,16'h002a,16'h0043,-16'h0132,-16'h0020,16'h0002,16'h0033,-16'h001f,16'h0043,16'h0065,-16'h00e2,16'h0024,16'h004a,-16'h0030,16'h000d,-16'h000a,16'h001e,-16'h00e1,-16'h000a,-16'h0035,-16'h0040,-16'h001a,-16'h0003,-16'h003c,-16'h001a,-16'h0003,-16'h0015,-16'h0003,16'h002f,-16'h0014,-16'h0032,-16'h0032,-16'h002b,16'h0007,-16'h0037,-16'h005a,-16'h0023,-16'h0001,-16'h0018,16'h00c1,16'h00c3,-16'h001d,-16'h0078,16'h0038,16'h004f,16'h0016,-16'h0105,-16'h007e,16'h0006,-16'h0017,16'h005a,16'h000a,16'h001b,-16'h002e,-16'h0002,-16'h000a,-16'h0043,16'h006f,16'h000b,16'h0033,-16'h0037,16'h0000,16'h0010,-16'h001b,-16'h0019,16'h0036,16'h0018,-16'h010d,-16'h0054,-16'h000c,16'h000f,-16'h002f,16'h002e,16'h0077,-16'h00be,16'h0030,16'h0054,-16'h0055,16'h004e,-16'h0017,-16'h0003,-16'h0033,16'h0002,16'h002e,-16'h0032,-16'h0011,16'h0016,-16'h0028,16'h000d,-16'h0002,-16'h0007,16'h0000,16'h003e,-16'h0019,-16'h001a,-16'h0056,-16'h0080,16'h0011,-16'h004f,-16'h00c0,-16'h0038,-16'h0013,16'h001c,16'h00a3,16'h00af,16'h0005,-16'h0055,16'h0040,16'h0067,16'h0043,-16'h00bb,-16'h00b9,-16'h0036,16'h0004,16'h0049,16'h0035,16'h002d,-16'h001d,16'h0019,-16'h0019,-16'h0051,16'h007b,-16'h0010,16'h004d,-16'h001f,-16'h009a,-16'h0022,-16'h0014,-16'h0014,16'h0024,16'h003a,-16'h00ce,-16'h0047,-16'h0019,16'h0007,-16'h0026,16'h0035,16'h005b,-16'h008a,16'h005f,16'h0066,-16'h0084,16'h002f,16'h0000,-16'h000e,16'h0066,-16'h0031,16'h0081,-16'h001b,-16'h0038,16'h0024,-16'h0012,-16'h0016,-16'h0013,16'h0027,16'h001a,16'h0029,-16'h0010,-16'h0009,-16'h0046,-16'h007c,16'h0008,-16'h0001,-16'h0108,-16'h0029,-16'h003a,16'h001e,16'h00b9,16'h007f,-16'h0009,-16'h0057,16'h003a,16'h008f,16'h0029,-16'h00aa,-16'h0090,-16'h0042,16'h0039,16'h0059,16'h003b,16'h001d,-16'h0045,-16'h0024,-16'h0006,-16'h0046,16'h0061,-16'h002c,16'h0043,-16'h001b,-16'h0088,16'h001d,-16'h0028,-16'h0004,16'h0029,16'h000f,-16'h0095,-16'h0059,-16'h005e,-16'h0031,-16'h004b,16'h004b,16'h004d,-16'h004b,16'h0050,16'h0039,-16'h00cd,16'h005a,16'h0030,16'h0005,16'h00ac,-16'h0020,16'h0077,16'h0010,-16'h0041,16'h005f,-16'h0026,-16'h0010,-16'h002f,16'h0012,-16'h0034,16'h0037,16'h0013,-16'h003b,-16'h0013,-16'h0032,16'h0030,-16'h0001,-16'h00c6,16'h000a,-16'h0006,16'h0027,16'h00ec,16'h003d,16'h0010,-16'h002f,16'h004f,16'h00d2,16'h0028,-16'h0060,-16'h0079,-16'h002e,16'h0057,16'h0053,16'h000f,16'h0038,-16'h0064,-16'h0035,-16'h002d,-16'h0019,16'h005f,-16'h001c,16'h003f,-16'h003d,-16'h0086,16'h0052,-16'h0045,-16'h0023,-16'h0013,16'h005a,-16'h0072,-16'h001a,-16'h0025,16'h0008,-16'h0061,-16'h0006,16'h005d,-16'h003e,16'h0003,-16'h000a,16'h0015,16'h0051,-16'h0018,16'h0032,16'h0038,16'h0046,-16'h0029,-16'h0032,16'h001e,-16'h0025,16'h0011,16'h000d,16'h0042,16'h002f,-16'h0004,16'h0079,16'h0009,-16'h001e,-16'h0017,16'h0012,16'h0004,-16'h0018,-16'h0027,-16'h0041,16'h0029,-16'h001e,-16'h0027,16'h0030,16'h0010,16'h003f,-16'h006d,16'h0018,16'h0007,16'h0064,-16'h0047,-16'h0014,16'h0019,-16'h0003,16'h001e,16'h0020,-16'h0010,-16'h0045,16'h0007,-16'h0025,16'h002d,16'h0056,16'h0047,16'h001e,-16'h0014,-16'h0026,16'h0021,16'h0030,16'h0024,16'h0062,-16'h0070,-16'h002b,-16'h0021,16'h0041,-16'h0054,16'h000d,16'h0043,-16'h0059,16'h0002,16'h0030,-16'h001f,16'h0063,-16'h001d,16'h0016,-16'h000f,16'h003d,16'h0006,-16'h0029,16'h000d,-16'h0019,16'h0003,-16'h0029,-16'h001c,-16'h0012,-16'h0022,16'h006f,-16'h0013,-16'h0009,-16'h001c,16'h0016,-16'h0025,-16'h0030,-16'h003a,-16'h000e,16'h0009,-16'h0008,-16'h0035,16'h000f,16'h0018,16'h0049,-16'h0068,-16'h0005,16'h003d,16'h0039,-16'h0057,-16'h0008,16'h000c,16'h001d,16'h002b,16'h0044,-16'h005a,-16'h0021,16'h0005,16'h000d,16'h003c,16'h0040,16'h002e,16'h0020,-16'h0003,-16'h0024,16'h000f,16'h0009,16'h0004,16'h0037,-16'h003f,-16'h0047,-16'h0045,16'h003d,-16'h0059,16'h0017,16'h0037,-16'h0062,16'h0015,16'h0033,-16'h0032,16'h0023,16'h0005,16'h006d,-16'h000d,16'h0050,-16'h0012,-16'h002a,16'h0028,16'h0028,16'h001f,-16'h00a8,-16'h0032,-16'h000d,16'h001d,16'h004a,-16'h0019,16'h0003,-16'h0014,16'h0004,-16'h0011,-16'h0034,-16'h0031,16'h0016,-16'h0013,16'h0007,-16'h002e,16'h000b,16'h000a,16'h004d,-16'h0066,-16'h0001,16'h0050,16'h0039,-16'h005c,-16'h0019,16'h001d,16'h002d,16'h0031,16'h0033,-16'h004b,-16'h004d,16'h0000,16'h0028,16'h0026,16'h0052,16'h003a,16'h0031,16'h0017,-16'h0020,-16'h002b,16'h0004,-16'h0023,16'h001f,-16'h0030,-16'h0011,-16'h0034,16'h002e,-16'h0031,16'h0016,16'h0034,-16'h0039,16'h000b,16'h001a,-16'h003e,16'h0023,-16'h000b,16'h0059,-16'h0015,16'h0034,-16'h002e,-16'h0010,16'h001d,16'h0047,16'h0029,-16'h00c2,-16'h0039,-16'h001f,16'h0014,16'h0061,-16'h0010,-16'h001c,16'h0004,16'h001f,16'h000d,16'h0003,-16'h003e,16'h0018,-16'h0012,-16'h000d,-16'h0022,-16'h000e,-16'h0002,16'h004d,-16'h0049,16'h000f,16'h0021,16'h003d,-16'h0081,-16'h0020,16'h0012,16'h0040,16'h004c,16'h0032,-16'h0063,-16'h002d,-16'h000b,16'h000a,16'h002c,16'h0060,16'h0051,16'h0035,16'h0023,-16'h0012,-16'h000c,-16'h000b,-16'h0046,16'h0031,-16'h0019,-16'h001e,-16'h002a,16'h0057,-16'h0022,-16'h0013,16'h002c,-16'h000f,16'h0002,-16'h0014,-16'h0022,16'h003f,-16'h0011,16'h0016,-16'h0028,16'h004e,-16'h0003,-16'h000f,16'h000f,16'h0019,16'h0010,-16'h0071,-16'h00b3,-16'h000f,16'h0027,16'h008c,16'h000f,-16'h0026,16'h0014,16'h0025,16'h0027,16'h000e,-16'h0047,16'h0003,-16'h002a,-16'h0027,-16'h0026,16'h0015,-16'h0001,16'h0053,-16'h001f,-16'h001d,16'h0022,16'h001b,-16'h009c,-16'h0016,16'h0017,16'h007a,16'h0053,16'h003e,-16'h006e,-16'h0045,16'h0001,-16'h000b,16'h0047,16'h0051,16'h0043,16'h0036,16'h0004,-16'h0030,-16'h004b,16'h0003,-16'h0071,16'h0032,16'h002d,16'h0000,-16'h0036,16'h004e,-16'h003b,-16'h0004,16'h003e,16'h0055,-16'h000c,-16'h0011,16'h0004,16'h003c,-16'h0016,-16'h004c,-16'h0009,16'h0059,-16'h001d,-16'h001f,-16'h0009,16'h002f,16'h000b,-16'h0053,-16'h010c,16'h0013,16'h0014,16'h00a5,16'h0016,-16'h0006,-16'h0004,16'h0017,16'h002a,-16'h0012,-16'h0036,-16'h0007,-16'h0012,-16'h001b,-16'h000c,16'h001c,-16'h001e,16'h0011,16'h0006,-16'h0003,-16'h001f,16'h0046,-16'h00c7,16'h0004,16'h0002,16'h0080,16'h0069,16'h004f,-16'h007b,-16'h0060,16'h000e,-16'h0002,16'h0032,16'h0029,16'h0018,16'h0019,-16'h001c,-16'h0009,-16'h0023,-16'h0024,-16'h004b,16'h0022,16'h003f,-16'h002e,-16'h003a,16'h005b,-16'h0009,16'h000b,16'h0033,16'h0063,-16'h000e,-16'h0021,16'h0018,16'h0022,-16'h0015,-16'h00e5,-16'h0014,16'h003a,-16'h0009,-16'h002a,16'h0000,-16'h0009,16'h0009,-16'h0046,-16'h0085,16'h0002,16'h000d,16'h00a0,16'h0012,-16'h0029,-16'h0029,16'h0026,16'h003a,-16'h0007,-16'h0018,-16'h0030,16'h003c,-16'h0024,-16'h003c,-16'h0002,-16'h001e,-16'h000e,-16'h000a,16'h0001,-16'h0015,16'h003a,-16'h00bd,16'h000b,16'h0025,16'h009f,16'h0048,16'h0067,-16'h004e,-16'h0089,16'h0058,-16'h0013,16'h0039,-16'h000e,16'h0015,16'h0006,-16'h0035,-16'h0015,-16'h0003,-16'h0024,-16'h0014,16'h0015,16'h0031,-16'h006f,-16'h002b,16'h004b,16'h000b,-16'h0011,16'h003f,16'h0072,-16'h0010,-16'h002d,16'h000f,-16'h0004,16'h0025,-16'h0091,-16'h001c,16'h004d,16'h0000,-16'h001c,16'h0011,16'h000a,-16'h0021,-16'h0081,16'h0020,16'h0034,16'h0006,16'h009c,-16'h0005,-16'h0024,-16'h0031,16'h0039,16'h005f,-16'h001b,-16'h0012,-16'h000d,16'h0071,-16'h004f,-16'h0033,16'h0009,-16'h0037,-16'h000d,-16'h000f,16'h0031,-16'h001c,16'h0035,-16'h0087,16'h0013,16'h0038,16'h00ad,-16'h0008,16'h0053,-16'h006c,-16'h00b4,16'h0039,-16'h0013,16'h003c,-16'h005e,16'h0013,-16'h0008,-16'h0010,-16'h0004,16'h002a,-16'h0027,-16'h0004,-16'h0017,16'h0000,-16'h006b,-16'h0001,16'h0058,16'h003e,-16'h0024,16'h004a,16'h0054,-16'h0016,-16'h0040,16'h0027,-16'h0002,16'h001e,16'h000e,-16'h0025,16'h0034,-16'h000b,16'h0002,-16'h0024,16'h0019,-16'h0014,-16'h006d,16'h0035,16'h0044,-16'h0002,16'h008f,-16'h0011,-16'h0008,-16'h003b,16'h0030,16'h0061,-16'h0023,-16'h0004,16'h0024,16'h0052,-16'h003f,-16'h0028,16'h0005,-16'h002a,-16'h0013,-16'h002b,16'h001d,-16'h0022,16'h0029,-16'h0065,16'h0011,16'h0038,16'h00b0,-16'h0070,16'h003a,-16'h0069,-16'h00d6,16'h0019,16'h000f,16'h0027,-16'h0078,-16'h0014,-16'h0029,-16'h0006,-16'h001a,16'h002b,-16'h0031,16'h001c,-16'h001b,16'h000c,-16'h004e,16'h0038,16'h0027,16'h0048,-16'h000f,16'h001c,16'h0058,-16'h0012,-16'h0041,16'h0002,-16'h001a,16'h0005,16'h009d,-16'h000f,16'h0035,-16'h000e,-16'h0015,-16'h001a,16'h001d,-16'h0015,-16'h0043,16'h0054,16'h0011,-16'h0043,16'h007f,-16'h0027,-16'h0023,-16'h001b,16'h002d,16'h0070,-16'h0050,-16'h001a,16'h001a,-16'h001c,-16'h0025,-16'h002d,-16'h000d,-16'h0044,16'h0009,-16'h0018,16'h002b,16'h0000,16'h0010,-16'h000e,16'h0008,16'h0036,16'h008b,-16'h0083,16'h002f,-16'h003a,-16'h00e5,16'h0006,16'h003a,16'h0018,-16'h0032,-16'h0028,-16'h0041,16'h0009,16'h0003,16'h004d,-16'h002f,16'h0031,-16'h0032,16'h0002,-16'h004d,16'h004a,16'h0060,16'h0055,-16'h0006,16'h0015,16'h0002,-16'h0001,-16'h0061,-16'h0021,-16'h0030,16'h001d,16'h0090,-16'h002d,16'h004f,16'h0022,-16'h002b,-16'h0016,16'h000b,-16'h002a,-16'h001a,16'h0063,16'h000c,-16'h0031,16'h004f,-16'h0022,-16'h0020,-16'h0015,16'h0017,16'h006b,-16'h007b,-16'h0016,-16'h0015,-16'h0094,16'h0019,-16'h003f,16'h0024,-16'h0026,-16'h0011,16'h000e,16'h0056,16'h0007,16'h0016,-16'h000a,16'h0004,16'h0038,16'h00a7,-16'h006a,16'h002f,16'h000c,-16'h00d0,16'h0037,16'h001e,16'h000a,16'h0017,-16'h0010,-16'h0032,16'h0023,-16'h0004,16'h005a,-16'h0041,16'h0049,-16'h0025,-16'h000f,-16'h0040,16'h0055,16'h0043,16'h0066,-16'h000f,16'h0005,16'h002e,16'h0002,-16'h0035,-16'h0018,-16'h0014,16'h0000,16'h005a,-16'h0026,16'h003a,-16'h000b,-16'h0011,16'h0000,16'h0013,16'h000a,16'h0006,16'h0055,16'h0010,16'h0010,16'h007f,-16'h0023,-16'h0010,-16'h0021,16'h0008,16'h0092,-16'h0073,-16'h001f,-16'h0011,-16'h00c6,16'h0053,-16'h0032,16'h0000,-16'h0049,-16'h0035,16'h0014,16'h0067,16'h0005,16'h0006,16'h000f,-16'h0015,16'h0052,16'h008c,-16'h0038,16'h002c,16'h002a,-16'h00c2,16'h0061,16'h000e,16'h0005,16'h003e,-16'h0005,-16'h001e,16'h0028,-16'h0005,16'h0063,-16'h0032,16'h004d,16'h0000,-16'h0048,-16'h0030,16'h0056,16'h004d,16'h0060,16'h0026,16'h002a,16'h0036,16'h0022,-16'h0003,-16'h004a,-16'h002d,-16'h001e,16'h001a,-16'h0035,16'h0060,-16'h002e,-16'h0024,16'h000d,16'h0006,16'h0031,16'h001b,16'h004b,-16'h0001,16'h0043,16'h0093,-16'h001f,-16'h0040,16'h001b,-16'h0022,16'h0066,-16'h0062,-16'h001a,16'h0000,-16'h005d,16'h0098,-16'h0032,-16'h0018,-16'h0056,16'h0003,-16'h002d,16'h0028,-16'h001e,-16'h001d,16'h001e,-16'h002f,16'h003c,16'h0074,-16'h0039,16'h0023,16'h002f,-16'h0094,16'h0041,16'h000f,16'h0000,16'h0076,16'h000a,-16'h002e,16'h0039,-16'h0008,16'h003e,-16'h0036,16'h0025,-16'h000e,-16'h003b,16'h000b,16'h006b,16'h005d,16'h006b,16'h0006,16'h0037,16'h0015,16'h001c,16'h001b,-16'h001c,-16'h0043,-16'h0035,-16'h0075,-16'h0036,16'h0046,-16'h0032,-16'h000c,-16'h002e,16'h002b,16'h005c,16'h0038,16'h0029,16'h0012,16'h006b,16'h0082,16'h0019,-16'h0041,16'h003d,-16'h0039,16'h0031,-16'h0029,-16'h0028,-16'h0013,-16'h001c,16'h0048,-16'h0003,-16'h000f,-16'h0042,-16'h0017,-16'h0025,-16'h0016,16'h0004,-16'h0027,16'h0004,-16'h0052,16'h0022,16'h005d,-16'h0046,16'h0024,16'h0036,-16'h007d,16'h0058,16'h0000,-16'h000b,16'h006d,16'h0004,-16'h002e,16'h0033,-16'h0010,16'h0040,-16'h0029,16'h0002,-16'h0009,-16'h001d,-16'h0014,16'h005a,16'h0058,16'h0046,16'h0009,16'h0040,-16'h0029,16'h0038,16'h0003,-16'h0005,-16'h004d,-16'h003f,-16'h00a0,-16'h002c,16'h002a,16'h0000,16'h0012,-16'h0038,16'h0036,16'h0079,-16'h0004,16'h0032,16'h0000,16'h0075,16'h008c,16'h000d,-16'h002a,16'h003b,-16'h0015,-16'h002e,16'h000d,-16'h0030,-16'h0029,16'h0000,-16'h00a6,16'h0002,16'h0010,-16'h003c,-16'h003f,-16'h0012,-16'h0029,-16'h0026,-16'h0018,16'h000e,-16'h004c,16'h004c,16'h005f,-16'h002a,16'h0018,16'h0048,-16'h0078,16'h0044,16'h0012,-16'h0013,16'h0034,16'h0052,-16'h0017,16'h0012,16'h0011,16'h0041,-16'h0037,16'h0008,16'h0008,-16'h004e,16'h0002,16'h0068,16'h0057,16'h0067,16'h0023,16'h0028,-16'h0029,16'h0040,16'h000c,16'h0008,-16'h001f,-16'h0053,-16'h0022,-16'h0009,16'h0033,16'h0020,16'h0016,-16'h0046,16'h0049,16'h006a,16'h0035,16'h0003,-16'h000a,16'h003f,16'h0082,16'h0023,-16'h0031,16'h0013,16'h0012,-16'h003d,16'h003a,-16'h0037,-16'h0042,16'h0025,-16'h011a,16'h0035,16'h002d,-16'h0054,-16'h005a,16'h000c,-16'h0019,-16'h0048,-16'h0016,16'h0003,-16'h002d,16'h003c,16'h006b,16'h0002,16'h001e,16'h004b,-16'h0055,16'h0045,16'h0023,-16'h0039,16'h0026,16'h003d,-16'h0023,-16'h0017,-16'h0017,16'h002b,-16'h0043,-16'h0038,16'h0013,-16'h001f,16'h000a,16'h003d,16'h0048,16'h0046,16'h0031,16'h004b,-16'h0045,16'h0037,16'h001d,16'h0020,-16'h0027,-16'h0064,16'h000e,16'h0014,16'h002b,16'h0020,-16'h0001,-16'h004d,16'h002e,16'h0046,16'h0022,-16'h0020,16'h001b,-16'h0010,16'h0047,16'h004e,-16'h0025,-16'h004f,16'h0042,-16'h0046,16'h0042,-16'h001e,-16'h004f,16'h0003,-16'h005d,16'h0044,16'h0046,-16'h0065,-16'h001d,16'h002a,-16'h0026,-16'h004f,-16'h0019,-16'h0011,-16'h001a,-16'h000d,16'h0075,16'h000b,16'h0007,16'h003c,-16'h0049,16'h003e,16'h004a,-16'h0058,-16'h0033,16'h004c,-16'h001b,-16'h000e,-16'h0003,16'h001d,-16'h005c,-16'h0052,16'h004a,-16'h001b,-16'h002b,16'h0045,16'h0031,16'h004f,16'h004f,16'h006a,-16'h0032,16'h0022,16'h000d,16'h0043,-16'h0011,-16'h005c,16'h0050,16'h0054,16'h002c,16'h0031,16'h0006,-16'h006a,16'h0021,-16'h000d,16'h003e,-16'h0055,16'h0017,-16'h0028,16'h0036,16'h005b,-16'h003e,-16'h0053,16'h004e,-16'h0058,16'h004a,-16'h0067,-16'h0049,-16'h0021,16'h004f,16'h0032,16'h003d,-16'h0071,-16'h000e,16'h0016,-16'h003d,-16'h0056,16'h0007,-16'h0005,16'h0002,-16'h0025,16'h0066,16'h0031,16'h0012,16'h0038,-16'h002a,16'h0018,16'h0051,-16'h0068,-16'h005b,16'h0076,-16'h002b,16'h0002,-16'h0017,16'h0019,-16'h0049,-16'h0036,16'h0056,-16'h0030,-16'h0018,16'h006b,16'h0031,16'h0020,16'h0044,16'h004f,-16'h0022,16'h0030,16'h0000,16'h0049,-16'h0017,-16'h0059,16'h0024,16'h0073,16'h0011,16'h0045,16'h0011,-16'h0059,16'h0026,-16'h007e,16'h0025,-16'h0042,16'h0008,-16'h000b,16'h0037,16'h0063,-16'h0047,-16'h0079,16'h0013,-16'h0044,16'h0026,-16'h003b,-16'h0016,-16'h0021,16'h004b,16'h003b,-16'h0024,-16'h0094,16'h0002,16'h002c,-16'h003c,-16'h005a,16'h0033,-16'h001a,16'h001d,-16'h0022,16'h0054,16'h004b,16'h0007,-16'h0001,-16'h002e,16'h000b,16'h0052,-16'h0038,-16'h0041,16'h0057,-16'h0017,16'h0019,-16'h003a,-16'h0005,-16'h0033,-16'h002c,16'h0043,-16'h0064,-16'h0033,16'h004a,16'h0063,16'h001c,16'h002a,16'h0037,16'h0007,16'h0067,16'h0001,16'h0028,16'h0011,-16'h0049,16'h0031,16'h0052,-16'h0001,16'h0015,16'h001a,-16'h003f,16'h0035,-16'h0182,16'h0000,-16'h001a,-16'h000e,-16'h0017,16'h005a,16'h002e,-16'h002e,-16'h0049,16'h0017,-16'h004f,-16'h000e,-16'h0024,16'h0045,16'h0004,16'h004b,16'h0069,-16'h00b6,-16'h006a,16'h0006,16'h0003,-16'h0018,-16'h0050,16'h0000,-16'h0035,16'h0031,-16'h0034,16'h0053,16'h0033,-16'h0013,-16'h0001,-16'h0029,16'h0019,16'h0037,-16'h002a,-16'h0035,16'h007d,-16'h0008,16'h0020,-16'h0001,16'h0005,-16'h0048,-16'h0010,16'h0038,-16'h00c7,-16'h000e,16'h0059,16'h005d,16'h0024,16'h0016,16'h0049,16'h0015,16'h0047,16'h0007,16'h003d,16'h0021,-16'h001d,16'h0007,-16'h0038,16'h0003,16'h0011,16'h000e,-16'h0035,16'h001b,-16'h01a2,-16'h0013,-16'h0030,-16'h0019,16'h000b,16'h004c,16'h0010,-16'h0039,16'h002a,16'h0027,-16'h001e,-16'h002c,-16'h000f,16'h006c,16'h0005,16'h0050,16'h0047,-16'h00c0,-16'h0067,-16'h0015,16'h0000,16'h0021,-16'h004e,-16'h0024,-16'h004c,16'h0000,-16'h004b,16'h003c,16'h004e,16'h0011,-16'h001d,-16'h001e,16'h0028,16'h0015,16'h0009,-16'h0020,16'h0076,16'h0013,16'h002d,-16'h0006,16'h0035,-16'h003a,-16'h0017,16'h000e,-16'h015a,-16'h0011,16'h004a,16'h003a,16'h0004,16'h0024,16'h005e,16'h0014,16'h0051,16'h0026,16'h0010,16'h001a,-16'h0004,-16'h0016,-16'h00e4,-16'h0003,-16'h0033,16'h0001,-16'h0004,-16'h0003,-16'h0108,-16'h0016,-16'h004b,-16'h000c,16'h0016,16'h0067,-16'h000e,-16'h003c,16'h0056,-16'h0009,-16'h001c,-16'h0045,-16'h0012,16'h0083,16'h0002,-16'h0008,16'h0046,-16'h0063,-16'h0066,-16'h0021,16'h000a,16'h003d,-16'h001a,16'h001f,-16'h0049,16'h0022,-16'h004b,16'h0044,16'h002a,16'h0020,-16'h001e,-16'h0004,16'h001b,-16'h0011,16'h0037,-16'h0002,16'h006e,16'h0004,16'h004d,16'h0018,16'h0028,-16'h0059,16'h0010,16'h0017,-16'h0168,-16'h0031,16'h0049,16'h0034,16'h0013,16'h0027,16'h0063,-16'h000c,16'h0059,16'h0007,16'h000f,16'h0000,-16'h001e,-16'h000c,-16'h01b4,-16'h004a,-16'h0073,-16'h0007,16'h0000,-16'h002d,-16'h009d,-16'h002f,-16'h002a,-16'h0023,16'h000c,16'h007d,-16'h004a,-16'h002f,16'h0061,-16'h0005,16'h0007,-16'h0035,16'h000a,16'h003d,16'h0000,-16'h007c,16'h005f,16'h0008,-16'h0072,-16'h0040,16'h0002,16'h0072,-16'h0006,-16'h0047,-16'h0067,16'h000c,-16'h003a,16'h003e,16'h0017,16'h0026,-16'h0035,16'h000a,-16'h0012,-16'h0098,16'h0058,16'h0027,16'h0040,16'h0000,16'h0058,16'h0006,16'h0008,-16'h004d,16'h002b,16'h0037,-16'h0156,-16'h006b,16'h007f,16'h003a,-16'h001d,16'h0041,16'h0077,-16'h0044,16'h0041,16'h0031,-16'h000e,16'h0017,-16'h000c,-16'h0024,-16'h017e,-16'h004f,-16'h0062,-16'h0042,16'h001a,-16'h0026,-16'h0069,-16'h000d,-16'h0013,-16'h0031,16'h0013,16'h0056,-16'h0054,-16'h0007,16'h001f,-16'h0032,16'h0026,-16'h002d,-16'h0015,16'h0000,16'h0009,-16'h00b4,16'h007f,16'h0072,-16'h0032,-16'h0030,16'h0039,16'h0072,16'h000b,-16'h009c,-16'h008b,16'h0004,-16'h001e,16'h0050,16'h0015,16'h0029,-16'h0028,16'h0021,-16'h0033,-16'h0095,16'h006e,16'h003b,16'h002e,-16'h001c,16'h002d,16'h001a,16'h0007,-16'h0043,16'h0020,16'h0035,-16'h0126,-16'h0086,16'h005d,16'h000f,-16'h001c,16'h004a,16'h007d,-16'h005c,16'h003c,16'h0031,-16'h0016,16'h0027,-16'h001d,16'h0000,-16'h00f7,-16'h0025,-16'h001a,-16'h0048,16'h000d,-16'h0009,-16'h003a,16'h0004,-16'h0023,-16'h0027,16'h0018,16'h0047,-16'h0075,-16'h0022,-16'h0049,-16'h0038,16'h001e,-16'h0027,-16'h003c,-16'h005c,-16'h000d,-16'h0039,16'h0084,16'h00d4,-16'h000d,-16'h0050,16'h002c,16'h0070,16'h0005,-16'h00b1,-16'h008e,16'h0011,-16'h0003,16'h0046,16'h0020,16'h0027,-16'h0009,16'h0015,-16'h002e,-16'h0060,16'h005b,16'h0015,16'h003f,-16'h0043,-16'h0048,16'h001a,-16'h0028,-16'h002b,16'h000d,16'h002c,-16'h00f7,-16'h00c5,16'h0035,16'h002e,-16'h002f,16'h002a,16'h005d,-16'h006e,16'h0053,16'h0057,-16'h003d,16'h0035,16'h0012,16'h0017,-16'h000d,-16'h002e,16'h003a,-16'h003f,-16'h0004,16'h0029,-16'h001e,-16'h001a,-16'h0032,16'h0003,16'h001b,16'h0039,-16'h0079,16'h0006,-16'h006e,-16'h00b4,16'h003d,-16'h0027,-16'h0082,-16'h006e,-16'h001d,16'h0033,16'h00a9,16'h008b,-16'h0009,-16'h005f,16'h0039,16'h0059,16'h0035,-16'h006c,-16'h0092,-16'h001d,16'h0027,16'h0034,16'h001d,16'h0031,-16'h0013,16'h000e,-16'h0019,-16'h002b,16'h0072,-16'h0010,16'h0039,-16'h004a,-16'h00a3,-16'h0008,-16'h0013,-16'h0036,16'h0028,16'h0046,-16'h00c8,-16'h0092,16'h0002,16'h0020,-16'h0037,16'h003f,16'h0060,-16'h0051,16'h0055,16'h0057,-16'h0070,16'h0011,16'h001d,-16'h0020,16'h0073,-16'h0048,16'h0084,-16'h0043,-16'h0027,16'h003b,-16'h002f,-16'h0041,-16'h003c,16'h0038,16'h001b,16'h0029,-16'h002f,-16'h0013,-16'h0027,-16'h00fb,16'h003a,-16'h0006,-16'h00e8,-16'h005d,-16'h0020,16'h0025,16'h00ac,16'h006a,-16'h0016,-16'h007d,16'h0069,16'h0095,16'h0048,-16'h0074,-16'h0092,-16'h0032,16'h0032,16'h0028,16'h0018,16'h0045,-16'h004b,-16'h0003,16'h0010,-16'h0032,16'h0071,16'h0003,16'h004f,-16'h002a,-16'h008a,16'h0004,-16'h0009,-16'h002c,16'h0031,16'h002f,-16'h0091,-16'h008c,-16'h0048,-16'h0015,-16'h0055,16'h003d,16'h0048,-16'h004f,16'h0062,16'h0013,-16'h00af,16'h0044,-16'h0001,16'h001f,16'h00b4,-16'h003c,16'h009c,-16'h001b,-16'h0036,16'h003c,-16'h001b,-16'h003a,-16'h0031,16'h004a,-16'h0016,16'h0032,-16'h000a,-16'h003c,-16'h0009,-16'h009f,16'h0049,-16'h0025,-16'h00f6,-16'h0028,16'h000f,16'h003c,16'h00d6,16'h0017,-16'h002d,-16'h004e,16'h005a,16'h00ce,16'h002a,-16'h0067,-16'h0093,-16'h001b,16'h0066,16'h003c,-16'h0012,16'h0029,-16'h0048,-16'h0013,-16'h0011,-16'h0032,16'h0069,16'h0009,16'h005c,-16'h0014,-16'h0041,16'h0045,-16'h003d,-16'h001f,-16'h0004,16'h0071,-16'h0053,-16'h0023,-16'h003d,-16'h0011,-16'h0042,-16'h000b,16'h0061,-16'h002c,-16'h0016,16'h000b,16'h0003,16'h009f,-16'h0047,16'h002e,16'h0023,16'h0054,-16'h000e,-16'h0031,16'h001c,16'h0011,16'h0045,16'h0016,16'h001b,16'h0014,-16'h0030,16'h0066,16'h0015,-16'h0001,-16'h0029,-16'h0013,-16'h0003,-16'h0014,-16'h001f,-16'h0022,16'h0037,-16'h001a,-16'h0035,16'h0023,-16'h000e,16'h0069,-16'h0065,16'h002f,16'h001b,16'h0050,-16'h003d,-16'h0012,16'h0023,-16'h003b,-16'h0002,16'h0057,16'h0001,-16'h0012,-16'h001b,-16'h0036,16'h001a,16'h0051,16'h0040,16'h0039,-16'h0026,16'h000a,-16'h0002,16'h0042,16'h0027,16'h0072,-16'h005c,-16'h002d,-16'h0033,16'h000a,-16'h006e,16'h0011,16'h0064,-16'h0053,16'h0022,16'h0009,-16'h000a,16'h0063,-16'h0034,16'h006c,-16'h000f,16'h0046,16'h0033,-16'h0026,16'h0044,-16'h0005,16'h0035,-16'h001d,-16'h0021,-16'h0007,-16'h0017,16'h002a,16'h0000,-16'h0008,-16'h001b,16'h0009,-16'h000b,-16'h0014,-16'h002f,16'h0005,-16'h0006,-16'h001d,-16'h0038,16'h001a,16'h000f,16'h0044,-16'h006a,16'h000b,16'h004d,16'h0052,-16'h0032,16'h000a,16'h002b,-16'h0031,16'h0016,16'h004f,-16'h003f,-16'h002c,-16'h000b,16'h0003,16'h000d,16'h0044,16'h0057,16'h0017,16'h0024,-16'h0033,-16'h0016,16'h001f,16'h0016,16'h0067,-16'h0021,-16'h0030,-16'h0031,16'h0008,-16'h004c,16'h0019,16'h004f,-16'h0044,16'h0000,16'h0015,-16'h005b,16'h004b,-16'h001d,16'h0074,-16'h001a,16'h0055,16'h0016,-16'h002a,16'h0079,16'h0015,16'h0030,-16'h0089,-16'h0035,-16'h001c,16'h0017,16'h0034,16'h0001,-16'h0015,-16'h001c,16'h000a,16'h0010,16'h0001,-16'h0024,16'h0010,-16'h0011,-16'h000a,-16'h0044,-16'h0009,-16'h0022,16'h0067,-16'h0054,16'h0009,16'h003f,16'h002a,-16'h0042,-16'h0020,16'h001c,-16'h0001,16'h002e,16'h003c,-16'h0059,-16'h0016,16'h0003,16'h0016,16'h0023,16'h0055,16'h0050,16'h001d,16'h002a,-16'h0038,-16'h0036,16'h0004,-16'h0054,16'h0060,-16'h000e,-16'h0009,-16'h0017,-16'h0004,-16'h0066,16'h003e,16'h004b,-16'h0019,16'h002c,16'h0024,-16'h004b,16'h004a,-16'h0014,16'h0045,-16'h002c,16'h004a,16'h001a,-16'h0027,16'h006a,16'h004e,16'h002d,-16'h008b,-16'h0060,-16'h000d,16'h0016,16'h003f,-16'h0015,-16'h0010,16'h0007,16'h0019,16'h000b,16'h0002,-16'h0046,-16'h0016,-16'h0025,-16'h0032,-16'h0041,16'h0000,-16'h0006,16'h0059,-16'h0021,16'h000e,16'h003e,16'h0046,-16'h0063,16'h0003,16'h002c,16'h004e,16'h0039,16'h0039,-16'h0044,-16'h003d,16'h0008,16'h0020,16'h0045,16'h0048,16'h005e,16'h0030,16'h001a,-16'h0007,-16'h0025,16'h000d,-16'h0063,16'h003d,-16'h0008,-16'h0019,16'h0003,-16'h000b,-16'h0047,16'h001a,16'h005c,16'h002c,16'h0019,-16'h0002,-16'h0033,16'h006d,-16'h000b,16'h0021,-16'h0027,16'h005a,16'h003c,-16'h0017,16'h0069,16'h002e,16'h0029,-16'h0078,-16'h00a1,-16'h001a,16'h0001,16'h0062,16'h0008,-16'h001f,16'h0012,-16'h0010,16'h001c,16'h001f,-16'h0037,16'h0010,-16'h0022,-16'h0018,-16'h002f,-16'h0004,-16'h000b,16'h0044,-16'h001f,-16'h0009,-16'h0005,16'h003d,-16'h0074,-16'h0004,16'h0028,16'h0043,16'h0054,16'h0036,-16'h005e,-16'h0038,-16'h001f,16'h0021,16'h0047,16'h005b,16'h0053,16'h001c,16'h0005,-16'h0004,-16'h0032,-16'h0002,-16'h007d,16'h003a,16'h0031,-16'h0008,-16'h000d,16'h0015,-16'h0049,-16'h0011,16'h0055,16'h0062,-16'h000a,-16'h0016,-16'h0017,16'h006d,-16'h0009,-16'h0043,-16'h002c,16'h0051,16'h001e,-16'h0018,16'h006a,16'h0009,16'h001e,-16'h004d,-16'h00b0,16'h0005,-16'h000a,16'h006c,16'h0015,16'h0003,-16'h002a,16'h000f,16'h0069,16'h0029,-16'h0023,16'h0002,-16'h001e,-16'h0013,-16'h0016,16'h0019,-16'h0008,16'h0038,16'h0002,-16'h0026,-16'h0027,16'h0037,-16'h0083,16'h0004,16'h0038,16'h006f,16'h0040,16'h0055,-16'h0052,-16'h0059,16'h0005,-16'h000b,16'h0011,16'h004a,16'h004e,-16'h0007,-16'h0011,-16'h0005,-16'h0044,-16'h000b,-16'h003e,16'h0043,16'h0026,-16'h001d,-16'h0003,16'h0012,-16'h0043,16'h0000,16'h0055,16'h0073,-16'h0030,-16'h0036,16'h0004,16'h0079,16'h0025,-16'h00a8,-16'h0015,16'h0050,16'h0025,-16'h001d,16'h0062,-16'h001a,-16'h0014,-16'h0070,-16'h003d,16'h0005,16'h0002,16'h0090,16'h000c,-16'h0020,-16'h0023,16'h0001,16'h0044,-16'h001a,-16'h000b,-16'h000b,16'h0038,-16'h003d,-16'h0022,-16'h0001,-16'h0034,16'h0020,-16'h0013,-16'h0014,-16'h006b,16'h0040,-16'h008c,16'h0006,16'h003e,16'h0086,16'h0054,16'h004f,-16'h0034,-16'h0098,16'h004a,16'h0005,16'h0016,-16'h001e,16'h002f,16'h0002,-16'h0013,-16'h0008,-16'h0020,-16'h0026,-16'h0004,16'h0026,16'h0009,-16'h007a,-16'h0039,16'h0015,-16'h0048,16'h0009,16'h0035,16'h0043,-16'h0013,-16'h002b,16'h0000,16'h003e,16'h0023,-16'h0049,-16'h0033,16'h006f,16'h0011,-16'h001b,16'h0054,-16'h0008,-16'h001a,-16'h0064,16'h0035,16'h0026,-16'h002e,16'h0095,-16'h0003,-16'h000f,-16'h001d,16'h0027,16'h004e,-16'h000b,-16'h000c,-16'h000b,16'h008c,-16'h0035,-16'h002e,16'h0013,-16'h0051,-16'h0014,-16'h0028,16'h000c,-16'h0076,16'h0031,-16'h0081,16'h001e,16'h001c,16'h008a,-16'h0006,16'h0053,-16'h0068,-16'h00c9,16'h0037,16'h0013,-16'h0029,-16'h0070,16'h0019,16'h0011,16'h001d,-16'h0013,-16'h0003,-16'h001f,16'h002a,16'h0027,16'h000b,-16'h006b,-16'h0012,16'h0010,-16'h0036,-16'h0017,16'h003a,16'h0045,-16'h002d,-16'h0023,-16'h000b,16'h000c,16'h0030,16'h0064,-16'h001b,16'h0047,16'h000d,16'h001d,16'h0037,16'h000d,-16'h002a,-16'h003f,16'h003a,-16'h0016,-16'h0052,16'h008e,-16'h003e,-16'h0003,-16'h0023,16'h003b,16'h0069,-16'h004d,-16'h000e,16'h000e,16'h0048,-16'h005e,-16'h0039,16'h0007,-16'h0026,-16'h0016,-16'h0011,16'h001e,-16'h0038,16'h000d,-16'h004a,16'h0027,16'h0044,16'h008b,-16'h005d,16'h0048,-16'h004e,-16'h0100,16'h0020,16'h0038,-16'h001b,-16'h0070,16'h000e,-16'h0016,-16'h0014,-16'h0005,16'h0004,-16'h0025,16'h005d,16'h0008,-16'h000e,-16'h005b,-16'h000c,16'h0042,-16'h0027,-16'h0023,16'h0027,16'h0010,-16'h0008,-16'h001b,-16'h0011,-16'h0035,16'h0034,16'h00af,-16'h0007,16'h0053,16'h000f,16'h0003,16'h0037,16'h0020,-16'h0024,-16'h001f,16'h0054,-16'h001c,-16'h0042,16'h0058,-16'h003f,-16'h000b,-16'h0026,16'h0031,16'h0057,-16'h00bc,-16'h0039,16'h0003,-16'h005d,-16'h0042,-16'h0026,16'h0025,-16'h0032,16'h0017,16'h0013,16'h0052,-16'h0024,16'h001c,-16'h000c,16'h0040,16'h0056,16'h00a6,-16'h0057,16'h005a,-16'h002c,-16'h0115,16'h002b,16'h0028,-16'h004d,-16'h000c,16'h000c,-16'h0019,16'h002a,16'h0010,16'h001e,-16'h001a,16'h003c,-16'h002b,-16'h0016,-16'h004b,-16'h0004,16'h0041,-16'h002a,-16'h001e,16'h001f,16'h000c,-16'h0005,-16'h0041,-16'h0020,-16'h0048,16'h003b,16'h007e,-16'h0023,16'h0041,16'h0007,16'h000d,16'h0033,16'h0006,-16'h002b,16'h0034,16'h0051,-16'h0027,16'h0014,16'h0062,-16'h0035,-16'h001d,-16'h002a,16'h0029,16'h0058,-16'h00ed,-16'h0032,16'h002a,-16'h00c2,16'h0031,-16'h003a,16'h001e,-16'h0036,-16'h000a,16'h000a,16'h004f,-16'h0009,16'h0011,-16'h000c,16'h005b,16'h0051,16'h0073,-16'h000c,16'h0069,16'h0004,-16'h010f,16'h002b,16'h0017,-16'h001d,16'h0035,16'h0002,-16'h0035,16'h0046,16'h000d,16'h0023,-16'h001e,16'h004d,-16'h002b,-16'h0037,-16'h004d,16'h0009,16'h0041,-16'h001e,-16'h001b,16'h0029,16'h001a,16'h0007,-16'h0009,-16'h004b,-16'h0004,16'h0032,16'h002c,-16'h002e,16'h0035,16'h0026,16'h001a,16'h002a,16'h0026,-16'h0002,16'h0041,16'h0043,-16'h0024,16'h0045,16'h006c,-16'h0033,-16'h0010,-16'h0007,16'h0015,16'h008f,-16'h006b,-16'h0025,16'h000c,-16'h00b8,16'h006c,-16'h0030,-16'h0019,-16'h003c,-16'h0004,16'h0009,16'h006a,16'h0014,-16'h0015,16'h001d,16'h0051,16'h0081,16'h0080,-16'h001e,16'h006c,16'h0007,-16'h00e4,16'h0051,16'h000e,-16'h0014,16'h0055,-16'h0001,-16'h002e,16'h003b,16'h001b,16'h0037,-16'h0013,16'h0046,-16'h002f,-16'h0047,-16'h003c,16'h0016,16'h0035,-16'h0006,-16'h002e,16'h0013,16'h002a,16'h0023,16'h0022,-16'h004c,-16'h002d,16'h0014,-16'h0039,-16'h0030,16'h0029,-16'h0021,16'h0008,16'h002d,16'h001b,16'h003e,16'h0042,16'h001f,-16'h001b,16'h005f,16'h005f,-16'h000c,-16'h0033,16'h0045,-16'h0007,16'h0043,-16'h002d,-16'h002e,16'h001a,-16'h004a,16'h0075,-16'h0028,-16'h0021,-16'h0026,16'h000b,-16'h0021,16'h0037,16'h0005,-16'h003b,16'h0022,16'h0033,16'h0057,16'h004d,-16'h0008,16'h007e,16'h0021,-16'h00d2,16'h006c,16'h0023,-16'h0018,16'h007e,16'h0012,-16'h0017,16'h003d,16'h0000,16'h0042,-16'h0037,16'h0036,-16'h002b,-16'h003d,-16'h0046,16'h000a,16'h0044,-16'h0030,-16'h0024,16'h0031,-16'h0021,16'h0021,16'h0069,-16'h0019,-16'h0045,16'h0000,-16'h008e,-16'h0049,16'h0025,-16'h0024,-16'h000a,16'h0016,16'h001b,16'h0059,16'h0044,16'h0002,-16'h0004,16'h008d,16'h0084,-16'h0003,-16'h002a,16'h0041,16'h0000,-16'h0009,-16'h0009,-16'h0046,16'h0018,-16'h0013,-16'h0028,-16'h0046,16'h000c,-16'h0013,16'h0013,-16'h0039,-16'h0019,-16'h0006,-16'h0013,-16'h0008,16'h0029,16'h005d,16'h0048,-16'h0029,16'h0051,16'h0056,-16'h00c2,16'h0058,16'h0015,16'h0002,16'h0074,16'h0013,-16'h0009,16'h003a,16'h0006,16'h0032,-16'h002f,16'h0031,-16'h003b,-16'h0056,-16'h003a,16'h000a,16'h0048,-16'h0029,-16'h0012,16'h0011,-16'h005b,16'h0048,16'h0037,-16'h0016,-16'h0039,16'h0005,-16'h0055,-16'h004b,16'h000f,-16'h0002,16'h000a,-16'h0002,16'h003d,16'h0058,16'h0025,-16'h0006,-16'h000f,16'h0065,16'h0084,16'h0022,-16'h0020,16'h0022,16'h0007,-16'h0050,16'h002c,-16'h0050,-16'h001e,16'h000a,-16'h00f0,-16'h0016,16'h0004,-16'h002c,-16'h000d,-16'h0018,-16'h0033,16'h0004,16'h001f,16'h0004,16'h0030,16'h0044,16'h0050,-16'h0011,16'h0049,16'h0037,-16'h00b4,16'h004d,16'h0034,16'h000f,16'h0033,16'h0041,-16'h0006,16'h0008,16'h0002,16'h003d,-16'h003c,16'h001d,16'h0016,-16'h002f,-16'h001c,16'h000a,16'h0061,-16'h0021,16'h000b,16'h002d,-16'h0042,16'h0020,16'h0010,-16'h0013,-16'h001e,16'h0006,-16'h001a,-16'h0011,-16'h0002,16'h000d,16'h0011,-16'h001c,16'h0035,16'h0044,16'h0031,-16'h0059,-16'h0019,16'h0036,16'h0069,16'h002b,-16'h0016,16'h000b,16'h0029,-16'h004b,16'h0056,-16'h0048,-16'h006f,16'h002f,-16'h00ff,16'h0013,16'h003e,-16'h0028,-16'h0007,-16'h000f,-16'h0034,-16'h0013,-16'h0014,-16'h0009,16'h0022,16'h0046,16'h0048,-16'h0008,16'h003d,16'h002a,-16'h0095,16'h0057,16'h004c,-16'h0041,16'h002a,16'h0025,-16'h0003,-16'h0009,-16'h0007,16'h0038,-16'h0040,16'h0006,-16'h0009,-16'h001d,-16'h003c,16'h0014,16'h004d,-16'h0023,16'h0051,16'h0039,-16'h004f,16'h0037,16'h0021,16'h000e,16'h0022,-16'h0021,16'h006a,16'h0023,-16'h0004,16'h0011,-16'h0004,-16'h0010,16'h0030,16'h0014,16'h0025,-16'h0096,-16'h000d,-16'h000e,16'h006d,16'h005b,-16'h0035,-16'h0023,16'h0020,-16'h0064,16'h003a,-16'h004c,-16'h0088,16'h002d,-16'h0076,16'h0017,16'h0023,-16'h0038,16'h0014,-16'h0004,-16'h000e,-16'h003a,-16'h000e,-16'h0014,16'h0036,16'h0014,16'h0054,16'h002c,16'h000e,16'h001c,-16'h006d,16'h0047,16'h007a,-16'h0037,-16'h002a,16'h0023,-16'h0041,-16'h0014,16'h0010,16'h0037,-16'h004d,-16'h001d,16'h0001,16'h0000,-16'h0058,-16'h0008,16'h003f,-16'h000a,16'h004a,16'h002d,-16'h0041,16'h0037,16'h003f,16'h0038,16'h0016,-16'h002a,16'h0055,16'h004e,16'h0017,16'h0024,16'h0005,-16'h0015,16'h001c,-16'h0036,16'h0033,-16'h009f,-16'h0016,-16'h0029,16'h0055,16'h005b,-16'h001e,-16'h001a,16'h0010,-16'h0058,16'h0024,-16'h0059,-16'h0077,-16'h0011,16'h005a,16'h0007,16'h0038,-16'h003e,16'h0051,16'h000c,-16'h0042,-16'h0045,-16'h0003,-16'h0021,16'h000f,16'h0011,16'h003b,16'h0034,16'h0009,16'h0028,-16'h005f,16'h0047,16'h0093,-16'h002a,-16'h005a,16'h0024,-16'h0040,16'h0013,-16'h0010,-16'h000a,-16'h0047,-16'h0017,16'h0017,-16'h0001,-16'h0078,16'h0007,16'h0039,16'h000b,16'h002b,16'h001b,-16'h0006,16'h0035,16'h0011,16'h003b,16'h0002,-16'h001d,16'h0048,16'h007d,16'h000c,16'h0026,16'h0011,-16'h0007,16'h004f,-16'h0062,-16'h000b,-16'h0059,-16'h001b,-16'h001b,16'h004d,16'h0047,-16'h0034,-16'h002f,16'h0013,-16'h0041,-16'h0009,-16'h003e,-16'h0029,16'h0006,16'h0065,16'h0015,-16'h002e,-16'h004e,16'h0048,16'h000d,-16'h0044,-16'h006a,16'h0000,-16'h0051,-16'h001d,-16'h0016,16'h0028,16'h0045,16'h0000,-16'h000f,-16'h0054,16'h002a,16'h008d,16'h0031,-16'h003b,16'h002f,-16'h004b,16'h0031,-16'h0027,-16'h0010,-16'h0048,16'h0015,16'h001b,16'h0042,-16'h0058,16'h0005,16'h0032,16'h0000,16'h001e,16'h002d,16'h0019,16'h002a,-16'h0003,16'h0028,16'h001e,-16'h001d,16'h0037,16'h0062,16'h0006,16'h001a,16'h0023,16'h0004,16'h002e,-16'h00fb,-16'h0005,-16'h0043,-16'h000d,-16'h0024,16'h0033,16'h0020,-16'h0051,-16'h001d,16'h002f,-16'h0005,-16'h0028,-16'h0044,16'h002b,-16'h0005,16'h004f,16'h0032,-16'h0094,-16'h003d,16'h0049,-16'h0021,-16'h0005,-16'h0078,-16'h0027,-16'h0064,-16'h0021,-16'h001a,16'h000b,16'h004e,-16'h001e,-16'h0016,-16'h0052,-16'h001c,16'h004c,16'h0040,-16'h001d,16'h003b,-16'h003f,16'h005a,-16'h001d,-16'h0023,-16'h003b,16'h0013,16'h0026,-16'h0003,-16'h006d,16'h0012,16'h004a,16'h000d,16'h0016,16'h002b,16'h0016,16'h003f,16'h001b,16'h0022,16'h001a,-16'h0028,16'h0015,-16'h001d,-16'h0042,-16'h0006,16'h0022,16'h001e,16'h0005,-16'h016a,-16'h001f,-16'h0029,-16'h000a,16'h0008,16'h0033,16'h0010,-16'h004f,16'h0028,16'h0039,16'h000c,-16'h005f,-16'h0012,16'h0070,16'h0015,16'h0070,16'h0010,-16'h0094,-16'h0037,16'h001f,-16'h002a,16'h0045,-16'h0071,-16'h0038,-16'h006a,16'h0001,-16'h0007,-16'h001e,16'h0078,-16'h0012,-16'h0015,-16'h003f,16'h0001,16'h0015,16'h0043,-16'h000b,16'h0048,-16'h0015,16'h0077,-16'h0004,-16'h0007,-16'h0048,-16'h000f,16'h0004,-16'h0052,-16'h0084,16'h0036,16'h0041,-16'h001a,16'h002b,16'h0049,16'h0019,16'h0038,16'h0030,-16'h0002,16'h0015,-16'h0028,16'h0022,-16'h00d8,-16'h004a,-16'h003e,16'h001e,16'h0018,-16'h000b,-16'h010e,-16'h0030,-16'h001b,-16'h0004,16'h0016,16'h004f,-16'h0017,-16'h0038,16'h0046,16'h002d,16'h000e,-16'h003a,-16'h0009,16'h0065,16'h001f,-16'h000d,16'h0004,-16'h0065,-16'h0030,16'h0019,-16'h0015,16'h0053,-16'h002b,16'h000b,-16'h0064,16'h0014,-16'h001b,-16'h000b,16'h0040,16'h0011,-16'h0051,-16'h003a,16'h0019,-16'h007c,16'h005a,-16'h0013,16'h0038,-16'h001c,16'h0090,16'h0022,16'h001a,-16'h0046,16'h000f,-16'h0008,-16'h00b3,-16'h0091,16'h0079,16'h0017,-16'h0039,16'h004d,16'h0048,16'h002c,16'h0049,16'h0013,16'h0025,-16'h0015,-16'h003d,16'h0008,-16'h0179,-16'h0045,-16'h0053,16'h0023,16'h0030,-16'h0034,-16'h00a4,-16'h0009,-16'h0012,-16'h000d,16'h000a,16'h0055,-16'h004f,-16'h0021,16'h0041,16'h0006,16'h000c,-16'h0019,-16'h0023,16'h002c,16'h002d,-16'h00ac,16'h0009,16'h0017,-16'h002d,16'h0013,-16'h0003,16'h004b,-16'h000f,-16'h000d,-16'h0055,-16'h001c,16'h0014,-16'h0004,16'h0028,16'h0023,-16'h0039,-16'h0008,-16'h0017,-16'h00af,16'h006f,-16'h0001,16'h0028,-16'h0001,16'h0033,16'h0025,16'h0039,-16'h0042,-16'h0017,16'h0027,-16'h00fb,-16'h009c,16'h0073,16'h0025,-16'h002f,16'h007d,16'h0085,16'h0003,16'h003c,16'h001e,-16'h0021,-16'h0001,-16'h0023,-16'h0002,-16'h0165,-16'h0037,-16'h0024,16'h0000,16'h0051,-16'h002b,-16'h0075,-16'h0015,-16'h001e,-16'h0021,16'h0007,16'h006f,-16'h00b1,-16'h001e,16'h0019,-16'h0005,-16'h0016,-16'h0016,-16'h001a,-16'h002b,-16'h0001,-16'h00b0,16'h000c,16'h007a,-16'h0023,16'h0009,16'h0027,16'h0064,-16'h0005,-16'h0055,-16'h006b,-16'h0010,16'h0011,16'h0025,-16'h0003,16'h0036,-16'h0022,-16'h0026,-16'h0039,-16'h0069,16'h007f,16'h0009,16'h0029,-16'h0023,-16'h000d,16'h000a,16'h002b,-16'h003a,16'h0003,16'h0020,-16'h00b1,-16'h00d3,16'h0090,16'h0000,-16'h0015,16'h0050,16'h007c,-16'h0022,16'h0047,16'h0033,-16'h0020,16'h002d,16'h0006,16'h0005,-16'h00f7,-16'h0025,-16'h000d,-16'h004b,16'h0036,-16'h000e,-16'h004c,-16'h0028,-16'h003c,-16'h0033,16'h000a,16'h004f,-16'h0109,16'h0002,-16'h001c,-16'h0053,-16'h0021,-16'h0009,-16'h0053,-16'h007e,16'h0018,-16'h0035,-16'h0001,16'h00ba,-16'h0016,-16'h002a,16'h0005,16'h0059,-16'h000d,-16'h0085,-16'h0072,-16'h000b,-16'h0002,-16'h0005,-16'h0007,16'h004d,16'h0003,-16'h001f,-16'h003a,-16'h004b,16'h004b,16'h0013,16'h003d,-16'h002e,-16'h0086,16'h0014,16'h000c,-16'h003f,-16'h0003,16'h0005,-16'h00a3,-16'h00d5,16'h0065,-16'h0006,-16'h0027,16'h002b,16'h0042,-16'h0055,16'h0043,16'h002b,-16'h0008,16'h0018,16'h001a,16'h0003,-16'h001b,-16'h0029,16'h004a,-16'h0055,16'h0029,16'h000c,-16'h003b,-16'h003b,-16'h0018,16'h000c,16'h0016,16'h0065,-16'h00e0,16'h0002,-16'h0049,-16'h0102,-16'h0006,-16'h000e,-16'h005f,-16'h00b6,16'h0009,16'h0044,16'h0042,16'h0093,16'h0010,-16'h0041,16'h0009,16'h0064,16'h000a,-16'h004a,-16'h006f,16'h0007,16'h0017,16'h0000,16'h001c,16'h0059,-16'h0013,16'h0002,-16'h0040,-16'h000c,16'h005b,16'h000f,16'h0026,-16'h003f,-16'h00bc,-16'h0009,-16'h0005,-16'h0015,16'h0007,16'h004b,-16'h007a,-16'h00cc,16'h0040,16'h0006,-16'h0048,16'h0049,16'h005a,-16'h0039,16'h003d,16'h0057,-16'h002b,16'h0014,16'h0024,-16'h003e,16'h006c,-16'h0049,16'h008c,-16'h0048,-16'h001d,16'h0025,-16'h0034,-16'h0060,-16'h004b,16'h0014,16'h0030,16'h0047,-16'h006b,-16'h0018,-16'h003e,-16'h0134,16'h0013,-16'h0015,-16'h00a8,-16'h00a9,-16'h0006,16'h003d,16'h008d,16'h0022,-16'h0009,-16'h0059,16'h006d,16'h0072,16'h0068,-16'h004d,-16'h0065,16'h0024,16'h004d,-16'h0003,16'h002f,16'h004c,-16'h001d,16'h0016,16'h0000,-16'h0049,16'h006f,16'h0004,16'h0039,-16'h0030,-16'h005f,-16'h0032,-16'h002d,-16'h0013,16'h0028,16'h0040,-16'h005d,-16'h00e0,-16'h0011,-16'h000a,-16'h0064,16'h002d,16'h0057,-16'h0016,16'h0062,16'h0038,-16'h0042,16'h0050,16'h0008,-16'h001d,16'h00b5,-16'h005a,16'h0066,-16'h0040,-16'h0027,16'h0060,16'h0000,-16'h005f,-16'h0046,16'h0046,-16'h0003,16'h003c,-16'h0009,-16'h003c,-16'h001e,-16'h00ba,16'h0036,-16'h000d,-16'h00d3,-16'h0062,16'h0015,16'h004e,16'h00b2,-16'h000e,-16'h0025,-16'h006e,16'h0078,16'h0098,16'h0062,-16'h0047,-16'h0069,16'h001f,16'h0088,16'h0028,16'h002d,16'h002e,-16'h0052,-16'h0014,-16'h0010,-16'h005c,16'h0039,16'h000a,16'h0067,-16'h0038,-16'h001a,16'h0016,-16'h005b,-16'h002a,-16'h0011,16'h0066,-16'h0043,-16'h0005,-16'h0050,-16'h003a,-16'h0050,-16'h000f,16'h0075,-16'h001c,-16'h0007,-16'h0007,16'h0016,16'h009f,-16'h0025,16'h003f,16'h0020,16'h0037,16'h0009,-16'h0011,-16'h000d,16'h0003,16'h0038,-16'h0001,-16'h000c,16'h0002,-16'h001c,16'h0018,-16'h000c,16'h0020,-16'h0024,16'h0006,16'h0023,-16'h0017,-16'h0007,-16'h002e,16'h003d,-16'h0005,-16'h0015,16'h0011,-16'h0010,16'h007d,-16'h003d,16'h0019,16'h004c,16'h0066,-16'h000a,-16'h003e,16'h001c,-16'h004a,16'h0005,16'h005a,-16'h0019,-16'h0021,-16'h0020,-16'h002a,16'h0012,16'h004f,16'h0061,16'h004f,-16'h0003,-16'h0032,16'h0029,16'h0040,-16'h0011,16'h009b,-16'h0011,-16'h0012,-16'h0033,-16'h0032,-16'h0044,16'h0007,16'h0052,-16'h0035,16'h001d,-16'h0006,-16'h0028,16'h008a,-16'h0018,16'h004c,16'h0001,16'h0042,16'h0029,-16'h0035,16'h002d,16'h0016,16'h0017,-16'h001a,-16'h0046,-16'h0010,-16'h0001,16'h000a,-16'h0012,-16'h000c,-16'h0021,-16'h0007,16'h0003,-16'h0002,-16'h0009,16'h0000,16'h0008,16'h0002,-16'h0041,16'h0004,16'h000b,16'h0064,-16'h005f,-16'h000a,16'h005d,16'h0052,-16'h0034,16'h000a,16'h002c,-16'h002a,16'h0013,16'h003e,-16'h001e,16'h000f,-16'h001c,16'h001c,-16'h001b,16'h0054,16'h0069,16'h0021,16'h0013,-16'h0025,16'h0000,16'h0048,-16'h000e,16'h0083,16'h0004,-16'h000b,-16'h001d,-16'h004d,-16'h0052,16'h0025,16'h0040,-16'h0026,16'h0024,-16'h0002,-16'h0062,16'h0080,-16'h001a,16'h0054,-16'h0026,16'h005c,16'h0016,-16'h002a,16'h0059,16'h0016,16'h0022,-16'h0062,-16'h0049,-16'h001f,16'h0001,16'h0019,-16'h0020,-16'h0010,-16'h0025,16'h000c,16'h0025,16'h0022,-16'h000c,16'h0017,-16'h001e,16'h0002,-16'h0027,-16'h0006,-16'h002d,16'h004e,-16'h005b,16'h0003,16'h0053,16'h0055,-16'h0017,-16'h0017,16'h0045,16'h0001,16'h001f,16'h003b,-16'h0049,-16'h0010,-16'h0011,16'h0009,16'h0034,16'h0069,16'h005c,16'h001e,16'h002c,-16'h0010,16'h0006,16'h002e,-16'h004d,16'h0058,-16'h0004,16'h0008,-16'h0027,-16'h006c,-16'h003d,16'h0026,16'h006c,16'h0006,16'h001c,-16'h000d,-16'h006c,16'h0061,-16'h0001,16'h002f,-16'h0021,16'h0041,16'h004f,-16'h0015,16'h008d,16'h0057,16'h0033,-16'h0089,-16'h0066,-16'h0018,16'h0024,16'h0025,-16'h000e,-16'h0023,-16'h0007,-16'h000a,16'h0011,16'h003b,-16'h003d,16'h0020,-16'h003d,-16'h000b,-16'h0068,-16'h001d,-16'h002c,16'h0068,-16'h000b,16'h0003,16'h0007,16'h0044,-16'h0025,-16'h0001,16'h0011,16'h0039,16'h0021,16'h0041,-16'h0021,-16'h0014,16'h0008,16'h0011,16'h0021,16'h0052,16'h0077,16'h0041,16'h0039,-16'h0008,-16'h000a,16'h0018,-16'h005b,16'h005c,16'h0006,-16'h0007,-16'h0009,-16'h006b,-16'h0064,16'h0014,16'h005f,16'h000c,16'h0020,-16'h0004,-16'h004b,16'h00a7,-16'h0006,16'h0000,-16'h0018,16'h005b,16'h004e,16'h0005,16'h00b1,16'h0038,16'h0022,-16'h009c,-16'h00a5,-16'h0015,-16'h0016,16'h0054,16'h0014,-16'h000b,-16'h0004,-16'h001a,16'h002e,16'h0027,-16'h002f,16'h0017,-16'h003f,-16'h0023,-16'h003b,-16'h000e,-16'h0023,16'h0058,16'h0011,16'h000a,-16'h0020,16'h003c,-16'h0016,16'h000e,16'h001d,16'h0036,16'h0028,16'h0035,-16'h005c,-16'h0036,16'h0001,-16'h0007,16'h000b,16'h005b,16'h0042,16'h0037,16'h000c,-16'h001b,16'h0000,16'h0015,-16'h004d,16'h0057,16'h0035,16'h0010,16'h0009,-16'h0078,-16'h003b,16'h000c,16'h0054,16'h0042,-16'h0008,-16'h002f,-16'h002f,16'h0087,-16'h000b,-16'h0072,-16'h0018,16'h004a,16'h004e,-16'h0008,16'h0084,-16'h0005,-16'h0001,-16'h0063,-16'h0073,-16'h0006,-16'h0034,16'h005d,-16'h0003,-16'h000d,16'h0001,-16'h0025,16'h0044,-16'h0005,-16'h0035,16'h0000,16'h0004,16'h000f,-16'h0027,-16'h0012,-16'h0022,16'h0037,-16'h001e,16'h0024,-16'h004f,16'h0026,-16'h0003,-16'h0014,16'h0021,16'h002f,16'h000a,16'h0052,-16'h0029,-16'h0045,16'h0015,-16'h0001,-16'h0019,16'h002d,16'h0012,-16'h0003,-16'h0002,-16'h0007,16'h000c,-16'h0003,-16'h0004,16'h004a,16'h001b,-16'h0014,16'h0012,-16'h0057,-16'h0043,16'h002e,16'h0045,16'h0031,-16'h0025,-16'h002e,-16'h001d,16'h0078,16'h0017,-16'h005f,-16'h000e,16'h004f,16'h003c,16'h0001,16'h0098,16'h0003,-16'h0005,-16'h004b,-16'h0001,16'h000a,-16'h0025,16'h0066,-16'h0010,-16'h001d,16'h000a,16'h0004,16'h004a,16'h0001,-16'h002a,-16'h0028,16'h004c,-16'h0030,-16'h002b,-16'h0001,-16'h002a,16'h0021,-16'h001e,16'h0008,-16'h008c,16'h0057,-16'h001b,16'h0007,16'h004d,16'h002d,16'h004b,16'h006b,-16'h0047,-16'h005e,16'h0031,16'h0013,-16'h0036,-16'h0030,16'h0026,16'h0006,16'h000d,16'h0001,16'h000b,-16'h000e,16'h0038,16'h0028,16'h000e,-16'h0059,-16'h001e,-16'h0073,-16'h0049,16'h0022,16'h003b,16'h002a,-16'h000d,-16'h0019,-16'h0012,16'h0012,16'h002a,-16'h000a,16'h000a,16'h004c,16'h0022,16'h000f,16'h00a2,-16'h0003,-16'h0010,-16'h004b,16'h0042,-16'h0013,-16'h0040,16'h0029,-16'h0024,-16'h0008,16'h0013,16'h0030,16'h003c,-16'h006a,-16'h0027,-16'h0010,16'h0077,-16'h002f,-16'h0031,-16'h000b,-16'h0047,16'h0000,-16'h0013,16'h001e,-16'h008b,16'h002a,-16'h0020,-16'h0007,16'h0032,16'h003d,16'h0018,16'h0063,-16'h002f,-16'h0048,16'h002a,-16'h0004,-16'h005c,-16'h005a,16'h0003,16'h002e,16'h0034,16'h0000,16'h0016,16'h0004,16'h0051,16'h003a,16'h000d,-16'h0063,-16'h003c,-16'h005a,-16'h005e,16'h0000,16'h0018,16'h0014,-16'h0004,-16'h000d,-16'h0032,16'h0011,16'h0018,16'h007f,16'h0003,16'h003c,16'h0023,16'h0016,16'h0063,16'h000c,-16'h0029,-16'h001d,16'h0025,-16'h0055,-16'h003e,16'h0027,-16'h0049,-16'h001d,-16'h0022,16'h0022,16'h003c,-16'h00ba,-16'h0051,16'h0010,16'h001d,-16'h004c,-16'h001b,16'h0000,-16'h0034,16'h000e,-16'h0020,16'h0054,-16'h0073,16'h000d,-16'h0013,-16'h000f,16'h0055,16'h0049,-16'h003b,16'h004b,-16'h0044,-16'h005b,16'h0019,16'h001f,-16'h007e,-16'h0063,16'h0012,-16'h0003,16'h002b,16'h0010,16'h000b,16'h0010,16'h0063,16'h001b,-16'h000b,-16'h007c,-16'h0044,-16'h0022,-16'h005a,-16'h0020,16'h002a,-16'h0010,-16'h0011,-16'h002f,-16'h0074,-16'h001e,16'h003b,16'h00a4,16'h0026,16'h002c,16'h0023,16'h001b,16'h007e,16'h0023,-16'h0026,16'h000d,16'h0049,-16'h005d,16'h0015,16'h0034,-16'h0066,-16'h003e,-16'h001e,16'h0015,16'h003e,-16'h00e9,-16'h0058,16'h0020,-16'h007e,-16'h0027,-16'h002b,16'h0011,-16'h0041,-16'h001f,16'h001a,16'h0053,-16'h003c,16'h0032,-16'h0034,16'h002e,16'h006d,16'h003e,-16'h0037,16'h006a,-16'h0003,-16'h0060,16'h0003,16'h0000,-16'h0078,16'h0015,-16'h0012,-16'h0018,16'h0048,16'h001a,16'h0003,-16'h0017,16'h004a,-16'h0022,-16'h001b,-16'h0040,-16'h0018,-16'h0006,-16'h004c,-16'h0008,16'h003d,-16'h000a,-16'h000b,-16'h001c,-16'h007f,-16'h0043,16'h001e,16'h0066,-16'h0017,16'h0025,16'h0033,16'h0011,16'h0094,16'h0026,-16'h0045,16'h0057,16'h0037,-16'h0047,16'h0055,16'h0030,-16'h004c,-16'h0015,-16'h001c,16'h0001,16'h0059,-16'h0097,-16'h005b,16'h0038,-16'h00cc,16'h0021,-16'h0023,16'h001b,-16'h0059,-16'h0008,-16'h0001,16'h003d,16'h000d,16'h0003,-16'h001b,16'h0025,16'h006e,16'h001b,-16'h0029,16'h0067,16'h000c,-16'h004a,16'h000e,-16'h0007,-16'h003e,16'h0043,-16'h001a,-16'h0018,16'h0043,16'h0023,16'h002f,-16'h000c,16'h0052,-16'h0036,-16'h003b,-16'h003a,-16'h0037,-16'h0004,-16'h004f,-16'h0028,16'h001e,16'h0019,16'h0000,16'h0020,-16'h007f,-16'h0047,16'h0011,16'h0009,-16'h0042,16'h0004,16'h0018,16'h000b,16'h0075,16'h0025,-16'h0012,16'h0045,16'h001d,-16'h0050,16'h008f,16'h002d,-16'h001b,-16'h0021,16'h0017,-16'h000f,16'h005d,-16'h004c,-16'h0070,16'h0033,-16'h00bb,16'h0066,-16'h001a,-16'h0010,-16'h0053,-16'h000d,-16'h0002,16'h002c,16'h002c,-16'h0015,16'h000a,16'h0049,16'h007c,16'h0032,-16'h001f,16'h0070,16'h0016,-16'h0065,16'h0037,16'h0007,-16'h0048,16'h0056,16'h0013,-16'h000f,16'h003b,16'h001d,16'h0043,16'h0006,16'h003a,-16'h0021,-16'h0019,-16'h0055,-16'h002b,16'h0002,-16'h007a,-16'h0018,16'h0016,16'h0011,16'h0023,16'h0034,-16'h0060,-16'h003b,16'h001b,-16'h005d,-16'h0061,16'h0009,-16'h0012,16'h0004,16'h0070,16'h001c,16'h0026,16'h0049,16'h0004,-16'h0033,16'h008f,16'h0024,-16'h0007,-16'h0040,16'h0045,-16'h0043,16'h0018,-16'h0022,-16'h006c,16'h000a,-16'h002d,16'h007c,-16'h0022,-16'h0031,-16'h003c,16'h0004,-16'h002f,16'h001b,16'h0030,-16'h0013,16'h000c,16'h0021,16'h005e,-16'h0004,16'h0003,16'h007b,16'h0053,-16'h0057,16'h0029,16'h000e,-16'h004e,16'h003f,16'h0000,-16'h001f,16'h0038,16'h001a,16'h0029,-16'h0010,16'h005b,-16'h002a,-16'h0038,-16'h003f,-16'h0038,-16'h0001,-16'h0084,16'h0015,16'h0029,-16'h0045,16'h0034,16'h0055,-16'h0057,-16'h003f,16'h0007,-16'h005d,-16'h0060,16'h0000,-16'h0032,-16'h0014,16'h007d,16'h0019,16'h003f,16'h0031,-16'h0014,-16'h002c,16'h005b,16'h0030,16'h0015,-16'h002d,16'h0059,-16'h001d,-16'h0032,16'h000e,-16'h0059,16'h0033,16'h0003,-16'h000e,-16'h0042,16'h0010,-16'h0058,16'h0032,-16'h002e,-16'h001a,16'h000f,16'h0009,-16'h0020,16'h0043,16'h003a,-16'h0009,-16'h000a,16'h006b,16'h0062,-16'h0065,16'h0043,16'h0017,-16'h0033,16'h004d,16'h0013,-16'h0022,16'h001b,-16'h001a,16'h0007,-16'h0024,16'h0048,-16'h001a,-16'h0034,-16'h004f,-16'h0045,16'h0005,-16'h008f,16'h000a,16'h0026,-16'h0035,16'h0019,16'h001c,-16'h005e,16'h0005,16'h0012,-16'h0010,-16'h0060,-16'h0008,16'h0013,-16'h000e,16'h004b,16'h0016,16'h0035,16'h0020,-16'h0036,-16'h0023,16'h0041,16'h003b,16'h0016,-16'h0032,16'h0050,-16'h002e,-16'h003b,16'h0010,-16'h006f,-16'h0018,16'h0002,-16'h00c6,-16'h0036,16'h0047,-16'h0040,16'h001c,-16'h001c,-16'h0030,16'h000b,-16'h0007,16'h000e,16'h003c,16'h0041,-16'h0012,-16'h0004,16'h0069,16'h003d,-16'h0046,16'h005a,16'h001b,-16'h0007,16'h002e,16'h0010,16'h001c,16'h0020,-16'h0002,16'h0021,-16'h003c,16'h007a,-16'h001f,-16'h0029,-16'h004b,-16'h0018,-16'h0006,-16'h0097,16'h0016,16'h0020,-16'h002a,16'h000d,-16'h0001,-16'h0014,16'h002b,16'h001f,16'h0023,-16'h000b,-16'h0015,16'h000f,16'h0000,16'h0034,16'h003d,16'h0019,16'h0038,-16'h0046,-16'h0038,16'h0000,16'h004e,16'h002c,-16'h002f,16'h004f,-16'h0008,-16'h004b,16'h001e,-16'h004d,-16'h0088,16'h0027,-16'h00d0,-16'h0008,16'h002b,-16'h001d,16'h0028,-16'h0036,-16'h0061,16'h0010,16'h0009,16'h000b,16'h0053,16'h0042,-16'h0007,16'h001c,16'h003d,16'h0012,-16'h005c,16'h004a,16'h005d,-16'h0001,16'h000a,16'h0018,16'h0011,16'h001a,-16'h0026,16'h000d,-16'h0055,16'h005a,16'h000f,16'h000e,-16'h003c,-16'h0021,-16'h000a,-16'h0048,16'h0062,16'h0035,-16'h002e,16'h0026,16'h0008,16'h000c,16'h0039,16'h0008,16'h005c,16'h0039,16'h0004,16'h0016,-16'h0013,16'h0038,16'h0027,16'h000a,16'h0022,-16'h0040,-16'h0039,-16'h0037,16'h004e,16'h0011,-16'h0051,16'h000f,16'h0002,-16'h0061,16'h0021,-16'h0058,-16'h00cb,16'h0002,-16'h001e,16'h0001,16'h0022,-16'h0029,-16'h0018,-16'h001a,-16'h0038,-16'h0031,16'h001d,16'h0021,16'h0035,16'h001f,-16'h000a,-16'h0002,16'h0025,-16'h0007,-16'h004c,16'h003c,16'h0064,-16'h0007,-16'h0047,16'h0001,-16'h0017,16'h0019,-16'h0022,-16'h0039,-16'h0056,16'h0020,-16'h000c,16'h0031,-16'h009a,-16'h0025,-16'h0002,-16'h0035,16'h0063,16'h0027,-16'h003c,16'h002a,16'h0005,16'h0020,16'h000e,16'h001a,16'h0043,16'h004a,-16'h000c,16'h0036,-16'h000f,16'h003e,16'h002b,-16'h001e,16'h0008,-16'h0048,-16'h0051,-16'h0023,16'h002f,16'h0009,-16'h003b,-16'h0016,16'h002c,-16'h003d,16'h0017,-16'h0039,-16'h00af,16'h0017,16'h002c,-16'h000e,16'h000f,-16'h0057,-16'h0004,-16'h001b,-16'h0032,-16'h0052,-16'h0012,-16'h0002,16'h0015,16'h000d,-16'h000d,16'h003c,16'h0032,-16'h000a,-16'h002e,16'h0024,16'h0083,16'h0016,-16'h003d,16'h0002,-16'h003b,16'h0022,-16'h0006,-16'h005d,-16'h003e,16'h0023,16'h001b,16'h003c,-16'h007a,-16'h0014,-16'h0011,-16'h003f,16'h0060,16'h0018,-16'h0013,16'h002b,16'h0021,16'h0034,16'h001d,-16'h0002,16'h003a,16'h005c,16'h0025,16'h0030,16'h000f,16'h005c,16'h0018,-16'h004a,-16'h0013,-16'h005a,-16'h0033,-16'h0030,16'h002e,16'h0018,-16'h002e,-16'h001d,16'h0039,-16'h0034,16'h0000,-16'h002e,-16'h0061,16'h0014,16'h005f,-16'h0012,-16'h0036,-16'h0037,16'h0015,-16'h0004,-16'h0005,-16'h0045,16'h0007,-16'h0039,-16'h0007,16'h0011,-16'h001a,16'h0028,16'h0026,16'h001e,-16'h004c,16'h0014,16'h0038,16'h005c,-16'h0048,16'h0006,-16'h004e,16'h0028,-16'h0017,-16'h0081,-16'h0047,16'h001c,16'h001f,16'h006f,-16'h007a,-16'h0018,16'h0004,-16'h0021,16'h004d,16'h003a,16'h0013,16'h003f,16'h0002,16'h0021,16'h0025,16'h0005,16'h002e,16'h005d,-16'h0004,16'h003a,-16'h0012,16'h0056,16'h000b,-16'h0095,-16'h0012,-16'h002b,-16'h003a,-16'h0036,16'h003e,-16'h0009,-16'h0059,-16'h0005,16'h0027,16'h0015,-16'h0013,-16'h0047,16'h0019,-16'h0015,16'h0068,-16'h0002,-16'h00a1,-16'h001c,16'h002b,-16'h0020,16'h0016,-16'h0053,16'h0007,-16'h007d,-16'h0014,16'h0009,16'h0004,16'h0038,16'h0001,-16'h0008,-16'h0036,16'h0000,16'h000c,16'h0067,-16'h0014,16'h0022,-16'h004b,16'h005a,-16'h0001,-16'h0082,-16'h003c,-16'h0001,-16'h001a,16'h0085,-16'h00ad,-16'h001a,-16'h000e,-16'h002f,16'h0023,16'h0049,-16'h0005,16'h0031,16'h0036,16'h0025,16'h0029,-16'h0008,16'h0017,16'h0000,-16'h0029,16'h000a,-16'h0024,16'h003d,-16'h003b,-16'h0131,-16'h004e,-16'h002f,-16'h0007,-16'h0008,16'h0028,-16'h0001,-16'h0048,16'h004b,16'h003e,16'h0021,-16'h004f,-16'h0043,16'h006d,16'h0037,16'h004d,16'h000f,-16'h0077,-16'h0031,16'h002b,-16'h002c,16'h005f,-16'h0055,16'h0016,-16'h0083,16'h0020,16'h0004,-16'h003e,16'h0037,16'h0001,16'h0000,-16'h0046,-16'h0016,-16'h0059,16'h0087,16'h0003,16'h001c,-16'h0069,16'h0079,-16'h000b,-16'h0063,-16'h005d,-16'h0039,16'h0012,16'h0054,-16'h00e7,16'h0011,-16'h0019,-16'h0025,16'h003b,16'h0041,-16'h0013,16'h0004,16'h0040,16'h001c,16'h002b,-16'h001f,16'h0007,-16'h00e5,-16'h004a,-16'h0018,-16'h0018,16'h0034,-16'h005d,-16'h011c,-16'h0030,-16'h0010,-16'h002e,16'h000f,16'h005c,-16'h000d,-16'h0036,16'h003b,16'h0034,-16'h000f,-16'h0036,-16'h002e,16'h0065,16'h0027,-16'h001c,-16'h0009,-16'h0051,-16'h000b,16'h001a,16'h0010,16'h0051,-16'h0050,16'h000e,-16'h0054,16'h0000,16'h001f,-16'h005f,16'h0046,16'h0011,16'h0001,-16'h001c,16'h0000,-16'h008e,16'h0092,16'h0003,-16'h0004,-16'h003c,16'h006c,-16'h0004,16'h0000,-16'h005f,-16'h0030,16'h0001,16'h001b,-16'h0101,16'h004a,-16'h0031,-16'h0053,16'h0053,16'h0046,-16'h000e,16'h0024,16'h001e,16'h001b,16'h000c,-16'h0039,16'h0009,-16'h0159,-16'h004a,-16'h002b,16'h0011,16'h0032,-16'h0041,-16'h00dd,-16'h0042,16'h0020,-16'h002e,16'h000a,16'h0046,-16'h00ae,-16'h0027,16'h0025,16'h001c,-16'h004a,-16'h001e,-16'h0046,16'h002e,16'h002a,-16'h00ca,16'h0017,-16'h0002,-16'h0004,16'h0042,16'h001e,16'h005e,-16'h0012,16'h001f,-16'h0041,16'h0019,16'h0024,-16'h004c,16'h0022,16'h0042,16'h0005,-16'h0009,-16'h0010,-16'h0093,16'h0070,16'h0020,-16'h001e,-16'h002b,16'h0004,16'h001b,16'h003a,-16'h005a,-16'h0043,16'h0020,-16'h001c,-16'h00d5,16'h0052,-16'h0036,-16'h002e,16'h006a,16'h0063,-16'h000e,16'h0023,16'h0025,-16'h000f,16'h0010,-16'h0014,16'h000b,-16'h015c,-16'h005c,-16'h002a,-16'h0008,16'h0056,-16'h0040,-16'h009e,-16'h003e,16'h002d,-16'h002b,16'h000e,16'h0043,-16'h0142,-16'h0010,16'h0021,-16'h0014,-16'h00a3,-16'h0003,-16'h0044,-16'h000f,16'h0014,-16'h00a1,16'h0002,16'h007b,-16'h001a,16'h001f,16'h0018,16'h0054,16'h000a,-16'h0030,-16'h0050,16'h001c,16'h0000,-16'h0036,-16'h0006,16'h0010,16'h000d,-16'h000d,-16'h002c,-16'h005c,16'h0049,-16'h0005,16'h0010,-16'h003c,-16'h0076,16'h0014,16'h0031,-16'h003b,-16'h002a,16'h0001,-16'h0023,-16'h00cb,16'h0053,-16'h0011,-16'h0030,16'h0047,16'h005e,-16'h001f,16'h0036,16'h001f,-16'h0008,16'h0013,16'h0002,16'h0004,-16'h00ea,-16'h001c,16'h000a,16'h0000,16'h0040,16'h0001,-16'h0077,-16'h004d,16'h0002,-16'h0027,-16'h0009,16'h0040,-16'h014c,-16'h002d,-16'h0022,-16'h0070,-16'h00ab,-16'h0003,-16'h0060,-16'h008d,16'h0020,-16'h0029,-16'h0012,16'h00ba,16'h0016,16'h0005,16'h0012,16'h0061,-16'h0018,-16'h005b,-16'h0047,16'h001e,16'h002c,-16'h0041,-16'h0018,16'h0055,-16'h0005,-16'h0008,-16'h001f,-16'h0028,16'h001c,16'h0009,16'h0027,-16'h0055,-16'h0068,16'h0028,16'h0013,-16'h0034,16'h000c,-16'h0007,-16'h0058,-16'h00c4,16'h0038,-16'h0029,16'h0001,16'h000e,16'h005c,-16'h000a,16'h0028,16'h0021,-16'h000b,16'h0047,16'h001d,16'h0007,-16'h0029,16'h0002,16'h0053,16'h0004,16'h003e,-16'h0010,-16'h0032,-16'h0019,-16'h0004,-16'h001f,16'h001b,16'h0050,-16'h00e5,-16'h0017,-16'h004e,-16'h0129,-16'h0069,16'h0020,-16'h0091,-16'h00ba,-16'h0016,16'h0040,16'h0030,16'h0073,16'h0004,-16'h0016,16'h0024,16'h0069,16'h001c,-16'h0040,-16'h0047,16'h001c,16'h0050,-16'h0045,16'h0004,16'h006a,-16'h001d,16'h0016,-16'h0041,-16'h0010,16'h001f,16'h000e,16'h0040,-16'h002b,-16'h0083,16'h0000,-16'h0004,-16'h0032,16'h0025,16'h0056,-16'h004c,-16'h00dc,16'h0040,-16'h0018,-16'h0047,16'h001b,16'h004c,16'h0015,16'h0016,16'h0029,-16'h000b,16'h0021,16'h001e,-16'h0011,16'h005e,-16'h004a,16'h0099,-16'h0047,16'h0003,16'h0020,-16'h001b,-16'h002f,-16'h0049,16'h0006,16'h0043,16'h006d,-16'h007e,-16'h0037,-16'h0049,-16'h0135,-16'h000b,-16'h0004,-16'h00b2,-16'h00e3,-16'h0027,16'h0054,16'h0057,16'h000b,-16'h0021,-16'h0043,16'h0068,16'h0058,16'h005a,-16'h0019,-16'h002b,16'h0035,16'h0065,-16'h0046,16'h0027,16'h0048,16'h0000,-16'h0023,-16'h0008,-16'h0038,16'h0021,16'h0000,16'h0063,-16'h0030,-16'h0054,-16'h002f,-16'h0031,-16'h0016,16'h0007,16'h007c,-16'h0070,-16'h00d6,16'h0035,-16'h0046,-16'h00a8,16'h002a,16'h005d,16'h0010,16'h004b,16'h0022,-16'h0040,16'h004e,-16'h000c,-16'h0003,16'h00ab,-16'h008e,16'h0054,-16'h0072,-16'h0025,16'h004d,-16'h0003,-16'h007c,-16'h0060,-16'h000e,16'h003b,16'h0066,-16'h001a,-16'h007f,-16'h0017,-16'h00e5,16'h000e,16'h0003,-16'h00cf,-16'h0074,-16'h000b,16'h004b,16'h008f,16'h000b,-16'h0048,-16'h006f,16'h008a,16'h00a0,16'h0072,-16'h003f,-16'h005d,16'h0035,16'h006b,-16'h0015,-16'h0001,-16'h0017,-16'h003b,-16'h0039,-16'h000c,-16'h0051,16'h0007,-16'h0005,16'h009f,-16'h003f,-16'h001d,16'h0001,-16'h0082,-16'h0036,-16'h0023,16'h0063,-16'h0020,16'h0000,-16'h0068,-16'h004b,-16'h0039,-16'h002e,16'h004b,-16'h003d,16'h0007,-16'h0028,16'h002c,16'h00d2,-16'h0024,16'h0023,16'h0041,16'h0032,16'h0004,-16'h0014,-16'h002d,-16'h0006,16'h000a,16'h0008,16'h0013,16'h0016,-16'h001c,-16'h002c,16'h0014,16'h0023,-16'h0012,16'h0019,16'h0011,-16'h0004,16'h0044,-16'h0031,16'h0024,-16'h0002,-16'h0027,-16'h000e,-16'h002b,16'h007a,-16'h003a,16'h000b,16'h0059,16'h005b,16'h000b,-16'h002d,16'h0002,-16'h0059,16'h0006,16'h002e,-16'h000f,-16'h0011,-16'h0015,-16'h006b,-16'h0029,16'h0053,16'h0044,16'h0033,-16'h0005,-16'h002f,16'h0026,16'h0039,16'h000d,16'h0071,-16'h0017,16'h0008,-16'h0053,-16'h006a,-16'h0021,16'h0001,16'h0068,-16'h0051,16'h0022,-16'h0021,-16'h0021,16'h00b2,-16'h001c,16'h0058,16'h0003,16'h0056,16'h000f,-16'h000b,-16'h0002,16'h000f,16'h001b,-16'h0037,-16'h0036,-16'h0011,16'h000a,-16'h000c,-16'h0010,-16'h0012,-16'h0025,16'h0013,16'h0041,16'h001c,16'h0041,-16'h001a,-16'h000d,16'h0017,-16'h0011,16'h0004,-16'h000a,16'h0063,-16'h001d,16'h0014,16'h0050,16'h003c,-16'h000e,-16'h0002,16'h0025,-16'h003b,-16'h0002,16'h003a,-16'h0023,16'h0015,-16'h0001,16'h0003,-16'h001a,16'h0045,16'h0034,16'h0043,16'h002b,-16'h0023,16'h0054,16'h003c,16'h0005,16'h0076,-16'h0010,16'h0008,-16'h003d,-16'h0085,-16'h0016,16'h001f,16'h0059,-16'h0027,16'h0025,-16'h002c,-16'h005a,16'h0071,-16'h0012,16'h0059,16'h0003,16'h0050,16'h001a,-16'h003a,16'h0028,16'h001b,16'h0023,-16'h007f,-16'h0052,-16'h0001,16'h002d,-16'h0019,16'h000e,-16'h000e,-16'h0025,16'h001e,16'h001b,16'h0036,16'h0019,16'h001c,-16'h002a,16'h0003,-16'h0046,16'h0001,-16'h004d,16'h0067,-16'h0026,-16'h0006,16'h005e,16'h0041,-16'h000d,16'h0007,-16'h000a,-16'h0002,-16'h0012,16'h0033,-16'h004d,16'h0017,16'h0008,16'h0004,-16'h0030,16'h0040,16'h0050,16'h0015,16'h0028,-16'h0026,16'h0043,16'h0047,-16'h000a,16'h0039,-16'h000e,16'h0011,16'h0000,-16'h00aa,-16'h001b,16'h0030,16'h0033,-16'h000e,16'h002b,-16'h0011,-16'h006d,16'h007b,-16'h0010,16'h000b,-16'h0008,16'h006f,16'h0023,-16'h0010,16'h0051,16'h0049,16'h004d,-16'h0081,-16'h0054,-16'h0013,16'h0019,-16'h0038,-16'h0002,-16'h001c,-16'h000d,-16'h0015,16'h0034,16'h000a,16'h0004,16'h0029,-16'h0037,16'h001b,-16'h0021,-16'h001a,-16'h0053,16'h006f,-16'h000e,16'h001c,16'h0019,16'h0059,16'h0007,16'h0019,16'h001a,16'h0021,16'h0009,16'h0036,-16'h0047,-16'h001d,16'h000e,16'h000a,-16'h0062,16'h004d,16'h0029,16'h001e,16'h0019,-16'h0010,16'h0039,16'h0048,-16'h0021,16'h0040,-16'h000a,-16'h0012,16'h000b,-16'h00cb,-16'h0009,-16'h0002,16'h0032,16'h0005,16'h0012,-16'h0010,-16'h006e,16'h0053,-16'h0015,-16'h0016,16'h0001,16'h003b,16'h001c,-16'h0004,16'h0062,16'h0047,16'h002d,-16'h009c,-16'h0083,16'h0010,16'h001c,16'h001d,-16'h000c,-16'h0019,16'h000e,-16'h0023,16'h0042,16'h002b,16'h0000,16'h0041,-16'h003e,16'h000c,-16'h0029,-16'h003f,-16'h006c,16'h0050,-16'h0012,16'h0034,-16'h0042,16'h003f,16'h0035,16'h002c,16'h002f,16'h0030,16'h002e,16'h004f,-16'h0022,-16'h000e,-16'h0014,-16'h0004,-16'h006a,16'h000d,16'h0049,16'h003b,16'h0009,16'h000a,16'h001c,16'h004f,-16'h0023,16'h0024,16'h0018,16'h0016,16'h0023,-16'h00d1,-16'h0029,16'h0024,16'h0027,16'h0014,16'h0009,-16'h0018,-16'h0053,16'h0054,16'h000c,-16'h0072,16'h0021,16'h003b,16'h0007,-16'h0008,16'h005c,16'h0020,16'h002c,-16'h0069,-16'h004b,16'h0000,-16'h0040,16'h002a,-16'h0003,-16'h001d,16'h0019,-16'h002a,16'h0031,16'h001b,-16'h0024,16'h001b,16'h0000,16'h001f,-16'h0027,16'h0006,-16'h0040,16'h003e,-16'h001c,16'h0031,-16'h0057,16'h0025,16'h0035,-16'h000f,16'h000e,16'h0013,16'h003c,16'h0048,-16'h0024,16'h0007,-16'h000e,-16'h0001,-16'h008d,-16'h000a,16'h0025,16'h001a,16'h002f,16'h0018,16'h003e,16'h003d,16'h0030,16'h0042,16'h002b,16'h000b,-16'h0010,-16'h00b6,-16'h0038,-16'h0004,16'h0039,16'h000b,-16'h0017,-16'h001e,-16'h0036,16'h0016,16'h0016,-16'h0065,16'h0030,16'h002f,-16'h0007,16'h0021,16'h008a,16'h0007,16'h0011,-16'h0058,16'h000c,-16'h0001,-16'h0035,16'h002b,-16'h0024,-16'h0032,16'h003c,-16'h0018,16'h0041,-16'h0040,-16'h003f,-16'h0015,16'h004b,16'h002b,-16'h002f,-16'h0007,-16'h0044,16'h0054,-16'h001f,16'h005c,-16'h008c,-16'h0001,16'h0029,-16'h0023,16'h0030,-16'h0007,16'h003d,16'h003c,-16'h0030,16'h0002,16'h0003,16'h0014,-16'h005a,-16'h0042,16'h0027,16'h001c,16'h003f,16'h0002,16'h0025,16'h0038,16'h0057,16'h002f,16'h0008,-16'h000b,-16'h0011,-16'h00a4,-16'h0043,16'h002d,16'h003e,16'h000f,-16'h0007,-16'h0033,-16'h0070,-16'h000e,16'h000f,16'h001d,16'h0031,16'h0031,16'h0013,16'h0009,16'h0060,-16'h000f,-16'h0020,-16'h0040,16'h003f,-16'h001b,-16'h0033,-16'h000a,-16'h0045,-16'h0029,-16'h0004,-16'h000e,16'h0031,-16'h0081,-16'h002e,16'h0008,16'h0050,-16'h0003,-16'h001a,16'h0016,-16'h002a,16'h000f,-16'h0020,16'h006f,-16'h0092,16'h0023,16'h0000,-16'h0032,16'h0037,-16'h002e,16'h0009,16'h0050,-16'h003a,16'h002d,-16'h0019,16'h0015,-16'h007c,-16'h0079,-16'h0006,16'h002f,16'h003e,-16'h0023,16'h0025,16'h0041,16'h0044,16'h0024,16'h0003,-16'h0025,-16'h0061,-16'h0076,-16'h0036,16'h0010,16'h0031,16'h0019,16'h0008,-16'h0018,-16'h0074,-16'h000f,-16'h0024,16'h0093,16'h005b,16'h0019,16'h0043,16'h0001,16'h0065,16'h0007,-16'h0037,-16'h0003,16'h002d,-16'h003f,-16'h0024,-16'h0012,-16'h004a,-16'h0025,-16'h0008,-16'h0012,16'h003b,-16'h00cf,-16'h0068,16'h0000,-16'h0008,-16'h001b,-16'h0020,-16'h001a,-16'h004e,16'h0011,-16'h0035,16'h004a,-16'h0073,16'h0044,16'h0006,-16'h000c,16'h0070,-16'h0031,-16'h002a,16'h0037,-16'h0015,16'h002f,-16'h004b,-16'h0006,-16'h0071,-16'h0063,16'h000b,16'h0016,16'h002c,16'h0010,16'h000d,16'h0043,16'h0062,16'h001b,-16'h000b,-16'h004c,-16'h0060,-16'h008b,-16'h0034,16'h001e,16'h004c,16'h000e,16'h001e,-16'h0054,-16'h0093,-16'h004d,-16'h0004,16'h008f,16'h004f,16'h0010,16'h0040,16'h0027,16'h0071,16'h001c,-16'h0067,16'h0042,16'h0026,-16'h003c,16'h0058,-16'h0034,-16'h0039,-16'h0030,-16'h0017,16'h000f,16'h001f,-16'h00cc,-16'h006a,16'h0038,-16'h0071,-16'h0018,-16'h000c,16'h002a,-16'h0049,16'h0000,16'h0004,16'h0025,-16'h004d,16'h0041,-16'h0007,16'h001c,16'h004e,-16'h004a,-16'h0022,16'h0067,16'h0024,16'h0023,-16'h0036,-16'h000a,-16'h0064,16'h0020,-16'h000c,-16'h0022,16'h0045,16'h002f,16'h000f,16'h0029,16'h0070,-16'h003c,-16'h0020,-16'h0049,-16'h003d,-16'h0052,-16'h0005,16'h001e,16'h0037,16'h001b,16'h0031,-16'h0035,-16'h009b,-16'h009e,-16'h0003,16'h0056,16'h0022,16'h0011,16'h0045,-16'h000a,16'h007d,16'h0032,-16'h0036,16'h0065,16'h0022,-16'h005c,16'h0085,-16'h001c,-16'h0035,-16'h001e,-16'h0019,16'h000e,16'h005b,-16'h0067,-16'h005d,16'h0051,-16'h00c6,16'h0045,-16'h001b,16'h001f,-16'h004c,16'h0021,16'h0018,16'h002c,-16'h002c,16'h0030,16'h0009,16'h001a,16'h004f,-16'h004f,-16'h0015,16'h0059,16'h000d,16'h003e,-16'h001b,-16'h0012,-16'h0035,16'h0046,-16'h0001,16'h0001,16'h0065,-16'h0004,16'h000d,16'h0039,16'h0032,-16'h0010,-16'h0020,-16'h0026,-16'h003c,-16'h0054,-16'h0011,16'h002d,16'h0039,16'h0043,16'h0016,-16'h000f,-16'h0094,-16'h0070,16'h0008,-16'h0041,-16'h0037,16'h0012,16'h002a,16'h0005,16'h0079,16'h004b,16'h000e,16'h0044,16'h001b,-16'h005c,16'h00b2,-16'h002e,-16'h002d,-16'h002c,16'h001b,-16'h0024,16'h0049,16'h000e,-16'h0095,16'h0039,-16'h00b2,16'h008b,16'h0004,-16'h001b,-16'h0049,16'h0034,-16'h0002,-16'h000b,16'h0010,16'h0034,16'h001e,16'h0027,16'h0020,-16'h006e,-16'h000a,16'h0066,16'h0003,16'h0046,16'h0018,16'h0020,-16'h003f,16'h0037,16'h001c,-16'h000b,16'h004b,-16'h000d,16'h001c,16'h0022,16'h0058,-16'h0010,16'h0007,-16'h0025,-16'h0058,-16'h0046,-16'h002f,16'h003a,16'h0067,16'h0009,16'h0046,-16'h0011,-16'h0070,-16'h0075,16'h0012,-16'h0057,-16'h0046,-16'h000f,16'h000c,-16'h0023,16'h00a1,16'h0044,16'h0026,16'h0030,-16'h000a,-16'h0040,16'h007b,-16'h0039,-16'h0028,-16'h0031,16'h003c,-16'h004c,-16'h001e,16'h0032,-16'h0071,16'h0045,-16'h0014,16'h008b,16'h0005,-16'h005e,-16'h0040,16'h005b,16'h0000,-16'h0020,16'h002b,16'h0014,16'h0019,16'h003a,16'h001f,-16'h0074,-16'h0005,16'h0055,16'h0040,16'h003b,16'h000f,16'h004a,-16'h0024,16'h0049,16'h000e,-16'h0004,16'h0025,-16'h000b,16'h000a,16'h0023,16'h005c,-16'h001a,16'h002f,-16'h0029,-16'h0064,-16'h0045,-16'h0065,16'h003b,16'h0057,-16'h003b,16'h000a,-16'h0002,-16'h0066,-16'h003e,16'h000b,-16'h0048,-16'h0042,-16'h0007,16'h0021,-16'h0031,16'h009c,16'h0025,16'h001b,16'h0036,-16'h0035,-16'h0032,16'h0080,-16'h0026,16'h0003,-16'h0030,16'h007c,-16'h004e,-16'h002f,16'h0051,-16'h004e,16'h0052,16'h0020,-16'h0023,-16'h0021,16'h000b,-16'h004a,16'h0037,-16'h0023,-16'h0004,16'h0035,16'h0018,-16'h001a,16'h001e,16'h0000,-16'h0098,16'h000a,16'h0064,16'h004f,16'h0013,16'h0010,16'h003d,-16'h001d,16'h0030,16'h0037,16'h0000,16'h0023,-16'h0007,-16'h0002,16'h0001,16'h007e,-16'h000e,16'h0001,-16'h0014,-16'h004e,-16'h004c,-16'h0095,16'h006b,16'h0046,-16'h0051,-16'h000c,-16'h002c,-16'h005a,16'h0023,16'h0002,16'h0022,-16'h0024,-16'h0018,16'h001d,-16'h002b,16'h0089,16'h0022,16'h001d,16'h0027,-16'h002c,-16'h003b,16'h0033,-16'h001f,16'h0017,-16'h0031,16'h0067,-16'h0024,-16'h0011,16'h004e,-16'h004e,-16'h0011,16'h0005,-16'h00a9,16'h0000,16'h003f,-16'h0069,16'h0030,-16'h0010,-16'h0017,16'h0031,16'h0019,-16'h0023,16'h0039,16'h000b,-16'h0088,-16'h0007,16'h0076,16'h0017,16'h0028,16'h002c,16'h0036,16'h0001,-16'h0002,16'h001b,16'h000a,16'h0027,-16'h0020,-16'h0022,-16'h001c,16'h0083,-16'h000a,16'h0020,-16'h001b,-16'h0025,-16'h0049,-16'h008b,16'h0060,16'h0035,-16'h0025,-16'h002b,-16'h003d,-16'h0002,16'h0044,16'h0014,16'h0055,16'h0009,-16'h0015,16'h0028,-16'h003b,16'h0064,16'h0022,-16'h0004,16'h001c,-16'h003d,-16'h002d,-16'h003a,-16'h000f,-16'h0006,-16'h0033,16'h005c,-16'h002b,-16'h001b,16'h0059,-16'h004d,-16'h0081,16'h0024,-16'h0080,16'h0015,16'h000b,-16'h003b,16'h0001,-16'h0028,-16'h0045,16'h0007,16'h0019,-16'h000c,16'h0092,16'h0002,-16'h005d,-16'h002a,16'h0065,16'h0002,16'h000a,16'h0011,16'h0059,16'h0026,16'h0014,16'h0013,16'h0012,16'h002b,-16'h0025,-16'h0043,-16'h0008,16'h006c,-16'h000e,16'h0031,-16'h0059,-16'h0051,-16'h003a,-16'h008c,16'h0097,16'h0043,-16'h0069,16'h0001,-16'h002e,16'h002b,16'h0034,16'h0000,16'h0046,16'h000c,-16'h0039,16'h0028,-16'h0034,16'h005f,16'h0037,16'h000d,16'h002f,-16'h004c,-16'h003e,-16'h0054,-16'h0003,16'h0010,-16'h0045,16'h0015,-16'h0002,-16'h0010,16'h0054,-16'h0037,-16'h00cd,16'h0030,-16'h0018,16'h0021,-16'h0009,-16'h001e,-16'h0016,-16'h0009,-16'h0024,-16'h0023,16'h0002,16'h0002,16'h0073,16'h0018,-16'h0058,-16'h0046,16'h0057,-16'h0009,16'h0004,16'h0005,16'h0024,16'h0041,-16'h0013,16'h0029,-16'h0005,16'h001a,-16'h0004,-16'h005d,-16'h0009,16'h0022,16'h000a,16'h0030,-16'h0077,-16'h0020,-16'h0048,-16'h007e,16'h0088,16'h0037,-16'h005a,16'h0034,16'h0017,16'h001a,16'h000f,16'h0018,16'h0036,16'h000c,16'h0009,16'h001f,-16'h004c,16'h0061,16'h002e,16'h0003,16'h0022,-16'h002e,-16'h0050,-16'h000c,-16'h0005,16'h0016,-16'h0021,16'h0000,16'h001f,16'h0024,16'h0015,-16'h0045,-16'h00b9,16'h0017,16'h0029,16'h0013,-16'h0001,-16'h0007,-16'h0053,-16'h0013,-16'h0004,-16'h0032,-16'h001d,16'h000e,16'h0037,16'h0025,-16'h0057,-16'h002e,16'h0066,16'h0017,16'h0002,16'h0020,-16'h000b,16'h0053,-16'h000a,16'h0002,-16'h0011,16'h004c,16'h0001,-16'h0066,-16'h002f,16'h0027,16'h0010,16'h0046,-16'h005d,-16'h000e,-16'h0064,-16'h0053,16'h0069,16'h003e,-16'h003f,16'h003a,16'h0027,16'h000f,16'h0002,-16'h0012,16'h0024,16'h004a,-16'h0001,16'h0049,-16'h0014,16'h003e,16'h002f,-16'h002e,-16'h0023,-16'h0024,-16'h0039,-16'h0032,16'h0010,16'h0013,-16'h003e,-16'h0026,16'h0035,16'h0023,16'h000f,-16'h0036,-16'h0045,16'h0026,16'h004e,-16'h0005,-16'h0015,-16'h0003,-16'h0045,-16'h0012,16'h0019,-16'h0021,16'h0012,-16'h003f,16'h0017,16'h0012,-16'h0055,-16'h0010,16'h0061,16'h002d,16'h0000,16'h0010,-16'h0051,16'h0047,-16'h001d,16'h0031,-16'h0017,16'h002d,-16'h000c,-16'h00ae,-16'h0029,-16'h0008,16'h0026,16'h0055,-16'h0096,-16'h002d,-16'h0041,-16'h003c,16'h006a,16'h004f,-16'h0022,16'h0061,16'h0035,16'h000b,16'h0003,16'h0004,16'h001a,16'h0045,16'h0002,16'h0028,-16'h002b,16'h0052,-16'h0015,-16'h005f,-16'h0007,-16'h0005,-16'h0052,-16'h003b,16'h0032,-16'h001d,-16'h004c,16'h0024,16'h0024,16'h0029,16'h0005,-16'h0034,16'h000f,16'h000a,16'h003b,-16'h000c,-16'h0040,-16'h0002,16'h0007,-16'h000a,16'h0027,-16'h0049,16'h000b,-16'h004f,-16'h0007,-16'h0002,-16'h0031,16'h0025,16'h0037,16'h0023,-16'h0019,16'h000d,-16'h0059,16'h0053,-16'h0011,16'h003b,-16'h0041,16'h0058,-16'h0007,-16'h00ab,-16'h0016,-16'h004c,16'h0010,16'h0046,-16'h00cd,-16'h0014,-16'h0050,-16'h003a,16'h004d,16'h0027,-16'h003d,16'h0019,16'h0051,16'h0029,16'h0029,-16'h0015,16'h0008,-16'h001c,-16'h0034,16'h002d,-16'h001e,16'h0036,-16'h0027,-16'h0105,-16'h002e,-16'h0024,-16'h0019,-16'h0027,16'h0047,-16'h0013,-16'h0035,16'h0041,16'h0051,16'h000b,-16'h0012,-16'h002b,16'h0070,16'h0007,16'h000d,-16'h000d,-16'h0058,16'h000e,-16'h0003,16'h0019,16'h003b,-16'h006c,16'h0031,-16'h0034,-16'h0005,16'h0015,-16'h0051,16'h0030,-16'h000b,16'h001a,-16'h0010,-16'h0009,-16'h005a,16'h0056,16'h001f,16'h0028,-16'h0025,16'h0049,-16'h0021,-16'h009b,-16'h0055,-16'h0098,-16'h0019,16'h0065,-16'h0117,-16'h0019,-16'h0065,-16'h0031,16'h0064,16'h002f,-16'h0053,16'h000f,16'h004d,16'h0026,16'h004a,-16'h002a,-16'h0002,-16'h00c1,-16'h003d,16'h001c,-16'h001a,16'h0026,-16'h0052,-16'h0147,-16'h005b,-16'h0018,-16'h002c,16'h002f,16'h0060,-16'h0061,-16'h001d,16'h0048,16'h0037,-16'h0045,-16'h0016,-16'h002c,16'h0064,-16'h000d,-16'h0061,-16'h0016,-16'h001a,16'h001c,16'h000b,16'h0017,16'h0068,-16'h0055,16'h004f,-16'h0038,-16'h0010,16'h000c,-16'h0085,16'h0026,16'h001c,16'h0022,16'h0000,-16'h0012,-16'h0071,16'h0068,16'h0025,16'h0014,-16'h0001,-16'h0012,16'h0015,-16'h0028,-16'h0056,-16'h00c4,-16'h000f,16'h0040,-16'h0109,16'h001e,-16'h0072,-16'h0049,16'h0061,16'h004f,-16'h002e,16'h0018,16'h0046,16'h0022,16'h0045,-16'h000d,-16'h0012,-16'h014d,-16'h007a,16'h0010,16'h000e,16'h001e,-16'h0044,-16'h00fe,-16'h006a,16'h0023,-16'h0026,16'h0014,16'h0048,-16'h00fb,-16'h0038,16'h002a,16'h0011,-16'h0063,16'h000a,-16'h0036,16'h0031,-16'h0023,-16'h00ba,-16'h001a,16'h0018,16'h0028,16'h0031,16'h002c,16'h0051,-16'h0011,16'h003a,-16'h0028,16'h002b,16'h0012,-16'h0078,16'h0031,16'h001e,16'h0007,-16'h0013,-16'h000f,-16'h0073,16'h0064,16'h002e,16'h0002,-16'h002d,-16'h0048,16'h000d,16'h0038,-16'h0029,-16'h007c,16'h0013,16'h0020,-16'h00b9,16'h0013,-16'h0090,-16'h0032,16'h0051,16'h005e,-16'h002f,16'h0020,16'h003d,16'h0016,16'h001c,-16'h0010,-16'h000a,-16'h0135,-16'h0058,-16'h0003,-16'h0002,16'h0035,-16'h0028,-16'h00c6,-16'h005c,16'h001b,-16'h0032,16'h001d,16'h0042,-16'h014e,-16'h0040,16'h0003,-16'h0003,-16'h00d8,16'h0017,-16'h002e,-16'h0036,-16'h0011,-16'h00a9,-16'h002c,16'h009f,16'h0025,16'h001a,16'h0022,16'h005e,16'h001e,16'h000d,-16'h002a,16'h0036,16'h003b,-16'h005b,-16'h0009,16'h0021,-16'h000c,16'h0006,-16'h000b,-16'h004e,16'h0030,16'h0011,16'h0010,-16'h0014,-16'h0077,-16'h0003,16'h0041,-16'h0038,-16'h001b,-16'h0001,16'h0016,-16'h00a2,16'h003b,-16'h0074,-16'h0033,16'h003e,16'h0061,-16'h000a,16'h0018,16'h0029,-16'h0007,16'h001e,-16'h0003,16'h001d,-16'h00f3,-16'h0010,-16'h0003,16'h0015,16'h0041,-16'h001a,-16'h0087,-16'h0088,16'h0013,-16'h0045,16'h0004,16'h0059,-16'h010d,-16'h0037,-16'h0026,-16'h0093,-16'h00fd,16'h001a,-16'h004c,-16'h00d1,16'h0015,-16'h001b,16'h0006,16'h009a,16'h000d,-16'h0011,16'h0019,16'h0035,-16'h0005,-16'h002f,-16'h0029,16'h0034,16'h0032,-16'h003f,-16'h000b,16'h003d,-16'h000d,16'h0010,16'h0024,-16'h0014,16'h000f,16'h0005,16'h0013,-16'h0019,-16'h0049,16'h000a,16'h004a,-16'h0041,-16'h0001,16'h0003,-16'h0028,-16'h00b2,16'h002a,-16'h002c,16'h0005,16'h001b,16'h0035,16'h0024,16'h0004,16'h0020,16'h0000,16'h0034,16'h0024,-16'h0025,-16'h0038,16'h000a,16'h004f,16'h0023,16'h002c,-16'h000b,-16'h004f,-16'h0033,-16'h000d,-16'h0060,16'h002e,16'h0084,-16'h00e4,-16'h0017,-16'h004f,-16'h016a,-16'h0095,16'h0029,-16'h0089,-16'h0100,-16'h0024,16'h0039,16'h002c,16'h005c,16'h0000,-16'h0004,16'h0028,16'h0052,16'h001a,-16'h0023,-16'h0008,16'h0010,16'h0054,-16'h003e,-16'h0007,16'h005e,-16'h001c,16'h0008,16'h0000,-16'h0018,16'h0019,-16'h000d,16'h0039,-16'h0028,-16'h0060,-16'h0016,16'h0009,-16'h001c,16'h0012,16'h0062,-16'h004d,-16'h00dd,16'h0020,-16'h003d,-16'h0017,16'h002d,16'h0045,16'h002f,-16'h0014,16'h003d,-16'h000b,-16'h0012,16'h0017,-16'h001c,16'h006f,-16'h004b,16'h0096,-16'h004a,16'h0027,-16'h000e,-16'h0014,-16'h0044,-16'h0030,-16'h0050,16'h0042,16'h006b,-16'h0076,-16'h002f,-16'h0059,-16'h0133,-16'h0048,16'h002d,-16'h00c2,-16'h00e8,-16'h0021,16'h0058,16'h0042,16'h0013,-16'h0013,-16'h0009,16'h005c,16'h0039,16'h0048,-16'h002d,-16'h0011,16'h005a,16'h003f,-16'h001c,-16'h0008,16'h003f,16'h0006,16'h0004,16'h0018,-16'h0015,-16'h000f,16'h001c,16'h0037,-16'h0014,-16'h0022,-16'h005a,-16'h0053,-16'h0011,16'h0012,16'h0097,-16'h005c,-16'h00dd,16'h0020,-16'h0042,-16'h006b,16'h001a,16'h002c,16'h000f,16'h0000,16'h0034,-16'h0048,16'h0047,-16'h0013,-16'h0006,16'h00a5,-16'h00a2,16'h0053,-16'h009e,-16'h0002,16'h0021,-16'h001a,-16'h0053,-16'h0066,-16'h0060,16'h004a,16'h0073,16'h000c,-16'h0093,-16'h0017,-16'h0100,-16'h0013,16'h000c,-16'h00cc,-16'h0092,16'h001f,16'h007b,16'h0067,-16'h002b,-16'h006a,-16'h0043,16'h009d,16'h0048,16'h0057,-16'h0022,-16'h0032,16'h0071,16'h0054,-16'h000a,-16'h000c,-16'h001d,-16'h0009,-16'h004b,16'h0005,-16'h0053,-16'h0045,16'h000a,16'h00a1,-16'h0035,-16'h002a,-16'h002d,-16'h00b8,-16'h0018,-16'h004c,16'h0058,-16'h001a,16'h0030,-16'h0074,-16'h0044,-16'h001f,-16'h001e,16'h0029,-16'h000c,-16'h0009,-16'h004c,16'h0026,16'h00c2,-16'h0012,16'h002f,16'h002a,16'h0038,-16'h0046,-16'h0001,-16'h0047,16'h001b,-16'h0020,-16'h0026,-16'h0008,16'h0015,-16'h0029,-16'h0063,-16'h0030,16'h0030,-16'h0029,16'h0047,16'h0034,16'h0013,16'h005b,16'h0008,16'h0030,-16'h0012,16'h0016,16'h0025,-16'h0053,16'h006d,-16'h0028,16'h000c,16'h002f,16'h006b,16'h0029,-16'h0046,16'h0023,-16'h005a,16'h0005,16'h002d,-16'h0007,-16'h0023,-16'h001a,-16'h006e,-16'h0078,16'h0061,16'h002b,16'h0041,16'h0014,-16'h001b,16'h0037,-16'h0006,-16'h003b,16'h0074,-16'h001f,16'h000e,-16'h004c,-16'h0058,-16'h0004,16'h000b,16'h0047,-16'h0027,16'h000e,-16'h0035,-16'h001a,16'h00ac,-16'h003b,16'h003d,16'h0003,16'h002d,-16'h002f,-16'h000a,-16'h003a,16'h002b,-16'h0028,-16'h002c,-16'h0055,16'h0015,16'h0011,-16'h0038,-16'h0032,16'h0003,-16'h000a,16'h001a,16'h0036,16'h0012,16'h0051,16'h0006,16'h0006,16'h0005,16'h000d,-16'h001a,-16'h0059,16'h0072,-16'h0025,16'h001a,16'h0059,16'h004e,-16'h0013,-16'h0007,16'h0021,-16'h002c,-16'h0013,16'h002b,-16'h0048,-16'h0001,-16'h000d,-16'h0048,-16'h0064,16'h0046,16'h0030,16'h002a,16'h0002,-16'h001c,16'h004b,16'h001f,-16'h0025,16'h0048,16'h0013,16'h0001,-16'h0055,-16'h0097,16'h0008,16'h0017,16'h0026,-16'h003b,16'h0018,-16'h004e,-16'h0050,16'h0092,-16'h001b,16'h0049,-16'h0013,16'h004a,-16'h0039,16'h0003,-16'h001c,16'h0017,16'h0019,-16'h0063,-16'h0029,-16'h0006,16'h0014,-16'h004b,-16'h002b,-16'h0004,-16'h0003,16'h0008,16'h0041,16'h0037,16'h004b,16'h0021,-16'h0023,16'h0000,-16'h0017,-16'h0001,-16'h007b,16'h0086,-16'h0013,-16'h0004,16'h0044,16'h002b,16'h001d,16'h0007,16'h0020,-16'h001c,16'h000c,16'h001b,-16'h0023,16'h0011,16'h0000,-16'h002c,-16'h0079,16'h0033,16'h001d,16'h002a,-16'h0008,-16'h0015,16'h0034,16'h0039,-16'h0024,16'h0044,-16'h0009,16'h000a,-16'h002e,-16'h009f,-16'h000b,16'h0012,16'h001d,-16'h0027,16'h0031,-16'h002c,-16'h0056,16'h0051,-16'h000e,16'h0034,16'h000e,16'h0047,-16'h0055,-16'h000b,-16'h002e,16'h002f,16'h0047,-16'h0057,-16'h0030,16'h0001,16'h001a,-16'h004a,-16'h0022,16'h0002,16'h001d,-16'h0018,16'h0038,16'h0003,16'h0017,16'h002e,-16'h001c,16'h0018,-16'h003e,-16'h001d,-16'h009e,16'h0056,16'h0011,16'h001f,16'h0031,16'h0054,16'h003f,16'h002b,16'h002b,-16'h001d,16'h002b,16'h0028,-16'h0023,16'h0000,16'h001d,-16'h0010,-16'h00cc,16'h0028,16'h000f,16'h002e,-16'h0011,-16'h0017,16'h005a,16'h0066,-16'h003b,16'h004d,16'h000a,16'h0016,-16'h001b,-16'h00bb,16'h0025,16'h0004,16'h0015,-16'h001e,16'h000c,-16'h0020,-16'h0066,16'h0023,-16'h000d,-16'h0048,-16'h0002,16'h0037,-16'h0087,-16'h000a,-16'h004b,16'h000e,16'h0042,-16'h0069,-16'h0056,-16'h0014,-16'h0010,-16'h004c,-16'h0008,-16'h0012,16'h0000,-16'h0038,16'h002f,16'h0009,16'h0022,16'h0044,-16'h0004,16'h001f,-16'h0018,-16'h0049,-16'h006d,16'h0057,16'h0001,16'h0043,-16'h000f,16'h002e,16'h0074,16'h005e,16'h0012,16'h000b,16'h0013,16'h0040,-16'h0021,16'h0004,-16'h000d,16'h001f,-16'h00b8,16'h0016,16'h0008,16'h0035,-16'h0018,16'h0003,16'h004d,16'h005d,16'h000b,16'h003d,16'h0046,-16'h0001,-16'h000b,-16'h00ef,16'h001c,-16'h0010,16'h0025,16'h0011,16'h0015,-16'h0001,-16'h0052,-16'h0026,-16'h0009,-16'h009f,16'h002e,16'h0029,-16'h0045,-16'h001d,-16'h0013,16'h0004,16'h0029,-16'h0061,-16'h001f,16'h0015,-16'h0076,-16'h0020,-16'h001e,-16'h000b,16'h0020,-16'h006d,16'h001b,-16'h0006,16'h0001,16'h0019,16'h002b,16'h004f,-16'h002a,-16'h0031,-16'h005c,16'h005a,-16'h0024,16'h0059,-16'h0051,16'h0000,16'h0071,16'h001b,-16'h000b,-16'h0028,16'h0020,16'h0044,-16'h001f,16'h0035,16'h0023,16'h0030,-16'h00ad,-16'h0017,-16'h0008,16'h000d,16'h0019,16'h0014,16'h003b,16'h0055,16'h0036,16'h0026,16'h0002,16'h0010,-16'h0003,-16'h00d9,-16'h000f,16'h0011,16'h0001,-16'h0012,16'h0014,-16'h0039,-16'h0058,-16'h005f,-16'h000f,-16'h0043,16'h0044,-16'h0001,-16'h0031,-16'h0026,16'h002f,-16'h0014,-16'h0005,-16'h0051,16'h0024,16'h0023,-16'h0073,16'h0001,-16'h0023,-16'h0020,16'h001b,-16'h0060,16'h0025,-16'h0071,16'h0002,-16'h000e,16'h0077,16'h0058,-16'h004e,-16'h0012,-16'h0059,16'h005b,-16'h0026,16'h0081,-16'h0064,16'h001a,16'h0077,-16'h0011,16'h0033,-16'h003d,16'h002e,16'h0018,-16'h0038,16'h0031,16'h002f,16'h0035,-16'h0080,-16'h003b,16'h0006,16'h0012,16'h001b,16'h001c,16'h0047,16'h0066,16'h004a,16'h001b,16'h000a,-16'h0006,-16'h0008,-16'h00c7,16'h0001,16'h0016,16'h001b,16'h0000,16'h000a,-16'h0054,-16'h0090,-16'h0070,-16'h000d,16'h0041,16'h0053,16'h0022,16'h000e,-16'h001e,16'h001e,-16'h000d,-16'h0052,-16'h003d,16'h003e,-16'h0038,-16'h0067,-16'h001b,-16'h000f,-16'h0032,16'h002b,-16'h003f,16'h0033,-16'h0097,-16'h001d,-16'h001c,16'h007f,16'h0025,-16'h0043,16'h001c,-16'h0053,16'h004f,-16'h0028,16'h0072,-16'h00a5,16'h0011,16'h0071,-16'h0026,16'h0062,-16'h0060,16'h0039,16'h000f,-16'h0013,16'h0048,-16'h0018,16'h0041,-16'h0091,-16'h00a0,16'h0000,16'h002d,16'h0038,16'h0002,16'h0024,16'h0071,16'h0048,16'h003f,-16'h0004,-16'h002f,-16'h000c,-16'h00c9,16'h0009,16'h0020,16'h001d,16'h0018,-16'h0014,-16'h004e,-16'h0080,-16'h0089,-16'h0036,16'h0091,16'h0038,16'h0010,16'h0032,-16'h0005,16'h001b,16'h0003,-16'h0075,16'h000b,16'h005b,-16'h0061,16'h0008,-16'h002b,-16'h0010,-16'h002a,16'h000d,-16'h0012,16'h0040,-16'h00a0,-16'h0019,16'h0006,16'h001e,-16'h000f,16'h0000,16'h0031,-16'h004b,16'h002a,-16'h0032,16'h002a,-16'h009f,16'h001d,16'h0049,-16'h0012,16'h004f,-16'h0080,16'h0006,16'h0011,16'h0006,16'h005b,-16'h002c,16'h0046,-16'h0085,-16'h008d,16'h0006,16'h0018,16'h001d,16'h004c,16'h000c,16'h0059,16'h002f,16'h0013,-16'h0011,-16'h0025,-16'h0027,-16'h009d,16'h001b,16'h0018,16'h0023,16'h001d,16'h000d,-16'h0062,-16'h007b,-16'h00b6,-16'h0047,16'h007a,16'h005f,16'h0010,16'h0018,16'h0018,16'h004c,16'h0016,-16'h004c,16'h004d,16'h0019,-16'h0057,16'h0067,-16'h0046,-16'h0010,-16'h003c,16'h0010,16'h001e,16'h0032,-16'h0039,-16'h0018,16'h001a,-16'h006e,-16'h0012,-16'h000b,16'h0028,-16'h0034,16'h0026,16'h0011,-16'h0043,-16'h00b7,16'h0024,16'h0046,16'h0022,16'h0022,-16'h0098,16'h0006,16'h0011,16'h0028,16'h0074,-16'h000a,16'h0053,-16'h004c,16'h0024,-16'h0001,16'h0015,16'h003f,16'h0024,-16'h002d,16'h007b,16'h001e,16'h0000,-16'h000c,-16'h002a,-16'h0032,-16'h0096,16'h0041,16'h0032,16'h003b,16'h001f,16'h0020,-16'h0035,-16'h006f,-16'h0100,-16'h001f,16'h0012,16'h0004,16'h0026,16'h0023,-16'h0005,16'h0045,16'h002b,-16'h0024,16'h004d,16'h0016,-16'h0067,16'h0084,-16'h003d,-16'h0024,-16'h003f,-16'h000f,16'h0025,16'h002d,16'h0028,-16'h0024,16'h0030,-16'h0083,16'h0054,16'h0019,16'h0022,-16'h0035,16'h004e,16'h0036,-16'h0041,-16'h0099,16'h0043,16'h0064,16'h0016,-16'h0002,-16'h0083,-16'h0002,16'h001d,16'h0008,16'h004b,16'h0008,16'h005f,-16'h002f,16'h0058,16'h000c,-16'h0001,16'h0025,-16'h0007,-16'h0002,16'h006a,16'h0009,-16'h0007,-16'h0007,-16'h0004,-16'h0014,-16'h0087,16'h0057,16'h003c,16'h0052,16'h0028,16'h003a,-16'h003a,-16'h0013,-16'h00d6,-16'h0003,-16'h0066,-16'h0062,16'h0005,16'h002c,-16'h000a,16'h0040,16'h0026,16'h001b,16'h003c,16'h001b,-16'h004b,16'h0084,-16'h0030,-16'h0027,-16'h002a,-16'h0016,16'h0015,16'h0034,16'h006b,-16'h004c,16'h005f,-16'h0070,16'h0077,16'h001e,-16'h004b,-16'h0035,16'h0069,16'h001c,-16'h0033,-16'h0063,16'h0045,16'h003a,16'h002a,-16'h000a,-16'h006c,16'h0017,16'h001d,16'h002a,16'h004c,16'h000c,16'h0066,-16'h002f,16'h0058,16'h0014,16'h0000,16'h0037,-16'h0003,16'h0006,16'h0083,16'h0040,16'h0018,16'h0012,-16'h002e,-16'h0007,-16'h007d,16'h0042,16'h0021,16'h004f,16'h0004,16'h000d,-16'h0050,-16'h000c,-16'h0053,-16'h0008,-16'h007a,-16'h0064,16'h0012,16'h0024,-16'h000b,16'h0055,16'h004a,16'h000a,16'h002f,-16'h000c,-16'h004b,16'h0061,-16'h0046,16'h0000,-16'h002e,-16'h000b,-16'h0034,-16'h0008,16'h0077,-16'h002e,16'h0030,16'h0001,16'h0043,16'h001e,-16'h006a,-16'h000e,16'h003f,16'h0038,-16'h0047,-16'h0028,16'h003d,16'h0038,16'h0026,-16'h0012,-16'h008c,16'h000d,16'h0026,16'h003f,16'h001c,-16'h0001,16'h0074,16'h0000,16'h0066,16'h002b,-16'h0002,16'h0028,16'h001c,16'h000b,16'h0096,16'h0030,16'h0016,16'h000d,-16'h0022,-16'h0011,-16'h0085,16'h0058,16'h0022,16'h004b,-16'h0022,-16'h000f,-16'h0033,-16'h0003,-16'h0014,16'h0018,-16'h002f,-16'h005e,-16'h0010,16'h001b,-16'h003a,16'h003c,16'h0021,16'h0003,16'h0036,-16'h0021,-16'h000a,16'h0034,-16'h0045,16'h0029,-16'h0052,16'h0054,-16'h0053,-16'h0020,16'h007f,-16'h001c,16'h002a,16'h0063,-16'h003b,-16'h0003,16'h000c,-16'h001e,16'h002f,16'h001c,-16'h0034,16'h000d,16'h005d,-16'h0012,16'h001b,-16'h004a,-16'h009e,16'h0008,16'h0026,16'h0015,16'h0021,-16'h0017,16'h005c,16'h000e,16'h004c,16'h0016,16'h0016,16'h0013,16'h0028,-16'h0016,16'h00a4,16'h004f,16'h0009,16'h0020,16'h0004,-16'h000b,-16'h0076,16'h0051,16'h0065,16'h0061,-16'h0012,-16'h0001,-16'h0037,16'h0008,16'h002e,16'h0028,16'h0025,-16'h0002,-16'h0012,16'h0008,-16'h0016,16'h0054,16'h0020,16'h0015,16'h0038,-16'h0032,-16'h000e,16'h0002,-16'h0013,16'h0033,-16'h0055,16'h0056,-16'h0047,-16'h0011,16'h008f,-16'h0016,-16'h002e,16'h004c,-16'h0098,16'h0004,16'h002c,-16'h0028,16'h0011,16'h0024,-16'h0064,16'h003d,16'h0020,16'h000c,16'h0031,-16'h0023,-16'h007c,16'h0008,16'h004f,16'h001e,16'h0022,-16'h0011,16'h005c,16'h0026,16'h0002,16'h0015,16'h0003,16'h0039,16'h0012,-16'h0034,16'h0087,16'h0077,16'h0022,16'h0016,-16'h0034,-16'h000b,-16'h006d,16'h0024,16'h0061,16'h003c,-16'h002a,16'h000f,-16'h0053,16'h0029,16'h0034,16'h0003,16'h006e,16'h003c,-16'h001d,16'h0028,-16'h0035,16'h0036,16'h001b,-16'h0014,16'h002f,-16'h0030,-16'h0026,-16'h003c,-16'h0022,16'h0024,-16'h004c,16'h0058,-16'h0033,-16'h0014,16'h0085,-16'h0011,-16'h0083,16'h002f,-16'h004a,16'h0010,16'h0006,-16'h0015,-16'h000a,16'h0026,-16'h0049,16'h004c,16'h0018,16'h0000,16'h0030,-16'h000e,-16'h0040,-16'h002c,16'h004f,16'h0012,16'h001e,16'h0000,16'h0009,16'h0038,-16'h001a,16'h002b,-16'h0006,16'h003f,16'h0038,-16'h003c,16'h007c,16'h004b,16'h0002,16'h0017,-16'h0068,-16'h0009,-16'h0064,-16'h0002,16'h005b,16'h004b,-16'h0025,-16'h000c,-16'h0028,16'h003c,16'h0031,16'h0007,16'h0054,16'h003d,-16'h0022,16'h000c,-16'h0040,16'h004a,16'h0020,16'h0008,16'h0031,-16'h002f,-16'h001c,-16'h0034,16'h0006,16'h0029,-16'h004f,16'h001d,16'h0009,16'h000c,16'h005c,-16'h0012,-16'h0090,16'h0037,16'h002f,16'h0022,16'h0004,-16'h0011,-16'h0024,16'h001a,-16'h0022,16'h0037,-16'h0006,16'h0013,16'h0048,16'h000d,-16'h004b,-16'h006c,16'h002d,16'h0000,16'h0007,16'h0039,-16'h0021,16'h0046,-16'h0035,16'h0011,-16'h0007,16'h0037,16'h002b,-16'h002d,16'h0061,16'h0035,16'h0011,16'h0037,-16'h0044,16'h000b,-16'h0069,-16'h0055,16'h0074,16'h0040,-16'h0054,16'h002e,16'h001e,16'h001b,16'h0002,16'h0001,16'h0042,16'h001e,-16'h0015,16'h000d,-16'h0052,16'h0030,16'h0020,-16'h000f,16'h0000,-16'h002f,-16'h0031,-16'h000c,-16'h0043,16'h0021,-16'h004e,-16'h0008,16'h0033,16'h0024,16'h004a,-16'h0008,-16'h00d3,16'h0012,16'h0037,16'h0006,16'h0003,-16'h0017,-16'h004e,-16'h0009,-16'h001f,16'h0047,16'h0000,16'h0008,16'h0020,16'h0034,-16'h0037,-16'h0057,16'h0037,16'h0006,-16'h000e,16'h0012,-16'h003f,16'h0041,-16'h0023,16'h0023,16'h0001,16'h003d,16'h0002,-16'h0040,16'h0049,16'h002f,16'h0006,16'h004a,-16'h004a,16'h0002,-16'h0068,-16'h0068,16'h004e,16'h0058,-16'h003f,16'h0062,16'h0017,-16'h000d,-16'h0038,-16'h000f,16'h0047,16'h003e,-16'h0028,16'h000c,-16'h005b,16'h0050,-16'h0003,16'h000d,16'h0005,-16'h000d,-16'h0045,-16'h000b,-16'h0015,16'h0007,-16'h0048,16'h0001,16'h0037,16'h004c,-16'h0003,-16'h0012,-16'h0017,16'h000a,16'h0057,16'h0002,-16'h001d,16'h0018,-16'h0057,-16'h000f,-16'h0024,-16'h000e,-16'h0007,-16'h0045,16'h0022,16'h001f,-16'h0047,-16'h0047,16'h0044,16'h0019,16'h000c,16'h001a,-16'h0046,16'h001a,16'h000f,16'h003c,-16'h0011,16'h003a,16'h0012,-16'h006a,16'h0057,-16'h001e,16'h0018,16'h0012,-16'h0045,16'h0002,-16'h005a,-16'h0060,16'h003f,16'h003a,-16'h0028,16'h005f,16'h003f,16'h0015,16'h0002,-16'h0019,16'h0023,16'h0017,-16'h0035,16'h001b,-16'h0053,16'h001f,-16'h0026,-16'h002e,-16'h000e,-16'h0004,-16'h004b,-16'h001c,16'h000e,-16'h0013,-16'h0044,16'h001d,16'h0042,16'h0046,-16'h002e,-16'h0006,16'h0021,-16'h0006,16'h003b,16'h0001,-16'h0025,16'h000e,-16'h0016,16'h001b,16'h0015,-16'h0023,16'h0024,-16'h0037,16'h0034,16'h0035,-16'h0025,-16'h0002,16'h0023,16'h0035,16'h0001,16'h000b,-16'h0052,16'h001c,16'h000c,16'h0041,16'h0007,16'h0033,16'h0011,-16'h0099,16'h0037,-16'h0055,16'h0003,16'h0023,-16'h008b,-16'h001d,-16'h0068,-16'h0074,16'h001d,16'h003f,-16'h0059,16'h004d,16'h0062,16'h0038,16'h0019,-16'h0035,-16'h0008,-16'h0044,-16'h0025,16'h0016,-16'h0055,16'h0024,-16'h0038,-16'h0098,-16'h0005,-16'h0032,-16'h0049,-16'h0006,16'h002f,16'h0006,-16'h0027,16'h003b,16'h0051,16'h002d,-16'h000c,-16'h0024,16'h0076,-16'h001e,-16'h0053,16'h0000,-16'h0036,16'h0019,-16'h0007,16'h0001,16'h002f,-16'h0033,16'h0020,-16'h003c,16'h001e,16'h0040,-16'h001b,16'h000d,16'h0022,16'h0024,16'h0001,16'h0013,-16'h004f,16'h0033,16'h001a,16'h0029,16'h000f,-16'h000e,-16'h000e,-16'h0076,16'h0012,-16'h0083,16'h0000,16'h0028,-16'h00bd,-16'h0006,-16'h0063,-16'h004b,16'h0041,16'h0033,-16'h004c,16'h0032,16'h0074,16'h003b,16'h0031,-16'h004b,-16'h0007,-16'h0092,-16'h005a,16'h001f,-16'h002a,16'h0008,-16'h0040,-16'h0111,-16'h0049,-16'h001d,-16'h0048,16'h0049,16'h0038,-16'h00b6,-16'h0036,16'h0035,16'h004e,-16'h0038,-16'h000e,-16'h000a,16'h0077,-16'h003d,-16'h0082,-16'h001c,-16'h002c,16'h000d,16'h0011,16'h0028,16'h0043,-16'h0043,16'h0024,-16'h0014,16'h0013,16'h0025,-16'h003c,16'h0012,16'h0020,16'h001d,16'h0000,16'h000d,-16'h0019,16'h004f,16'h000d,16'h0034,16'h0022,-16'h0057,-16'h0022,-16'h000e,16'h0014,-16'h00be,16'h0018,16'h0016,-16'h00ee,-16'h001a,-16'h0079,-16'h0028,16'h003c,16'h0029,-16'h001e,16'h001e,16'h0049,16'h004d,16'h002b,-16'h000d,16'h0007,-16'h00e1,-16'h006f,16'h0021,-16'h0004,-16'h0008,-16'h0028,-16'h013b,-16'h005e,16'h0006,-16'h0003,16'h0050,16'h0021,-16'h018f,-16'h004c,16'h0011,16'h0039,-16'h0062,16'h0015,16'h0006,16'h001e,-16'h0035,-16'h00c5,-16'h001a,16'h001a,16'h0025,16'h0024,16'h0007,16'h0046,-16'h0017,16'h0029,-16'h001a,16'h0038,16'h0024,-16'h0041,16'h0026,16'h0035,16'h0019,16'h000d,16'h0016,-16'h003d,16'h004c,16'h001f,16'h002f,-16'h0004,-16'h006e,16'h0008,16'h0034,16'h0012,-16'h00c5,-16'h0015,16'h002a,-16'h00c0,16'h0016,-16'h0092,-16'h0016,16'h0029,16'h0052,-16'h0013,16'h0035,16'h003c,16'h0022,16'h0016,-16'h0026,-16'h0004,-16'h011a,-16'h006f,16'h000a,-16'h0002,16'h0003,-16'h002d,-16'h00f1,-16'h0069,16'h0058,-16'h002b,16'h000e,16'h0014,-16'h0148,-16'h0042,16'h0013,16'h001b,-16'h00da,16'h0048,16'h0008,-16'h0060,-16'h000c,-16'h008d,-16'h002d,16'h006d,16'h004c,16'h0001,16'h001e,16'h000d,16'h0019,16'h001e,-16'h001a,16'h0038,16'h002d,-16'h0061,-16'h0005,16'h0038,-16'h0002,16'h0007,16'h0007,-16'h0025,16'h005a,16'h0037,16'h000e,-16'h001a,-16'h0042,-16'h000b,16'h0049,16'h003f,-16'h0053,16'h0007,16'h000f,-16'h00a5,16'h0026,-16'h0064,-16'h000d,16'h0016,16'h0037,-16'h0002,16'h0003,16'h0037,16'h0037,16'h0013,-16'h0007,16'h0024,-16'h00f0,-16'h0025,16'h000b,-16'h0010,16'h0034,16'h0000,-16'h009b,-16'h0057,16'h0031,-16'h003f,-16'h001b,16'h0028,-16'h00bf,-16'h003d,-16'h000d,-16'h00ab,-16'h00da,16'h0052,-16'h0004,-16'h0118,-16'h0016,16'h0016,-16'h0014,16'h0075,16'h000e,-16'h0010,16'h0033,16'h0020,16'h001d,-16'h0018,-16'h0010,16'h0025,16'h0058,-16'h0022,-16'h000f,16'h0042,-16'h0007,16'h0027,16'h001c,16'h0002,16'h0019,16'h000e,16'h0026,16'h0008,-16'h004f,16'h001d,16'h0050,16'h002b,-16'h0008,16'h0033,-16'h000c,-16'h00bf,16'h0024,-16'h003c,16'h0035,16'h002b,16'h002d,16'h0021,-16'h0030,16'h0026,16'h0026,16'h0013,16'h0003,-16'h0015,-16'h0054,-16'h0012,16'h003e,-16'h0021,16'h002b,-16'h0019,-16'h0066,-16'h0023,16'h0000,-16'h0075,16'h0017,16'h004b,-16'h00c6,-16'h0033,-16'h0031,-16'h0180,-16'h0097,16'h002d,-16'h001e,-16'h0153,-16'h0015,16'h0057,16'h0013,16'h002e,16'h000a,16'h002f,16'h0029,16'h003a,16'h0051,16'h000b,16'h0001,16'h0038,16'h0054,-16'h0011,16'h0002,16'h0067,-16'h0004,16'h0021,16'h0019,-16'h0017,16'h000d,-16'h0010,16'h000a,-16'h0002,-16'h0039,-16'h0016,16'h0004,16'h0021,16'h0029,16'h0051,-16'h0042,-16'h00a2,16'h004a,-16'h003f,-16'h0008,16'h0013,-16'h000d,16'h0041,-16'h0043,16'h0036,16'h002a,-16'h0025,16'h002c,16'h0010,16'h0069,-16'h0041,16'h0067,-16'h0071,16'h002b,-16'h0055,-16'h001b,-16'h004e,-16'h0032,-16'h00a8,16'h001f,16'h0062,-16'h006f,-16'h002c,-16'h0019,-16'h015b,-16'h003b,16'h0031,-16'h0059,-16'h00f9,-16'h0012,16'h0071,16'h0008,16'h0007,-16'h0034,16'h004e,16'h0057,16'h001f,16'h0072,16'h0003,16'h0012,16'h005f,16'h0059,-16'h002c,16'h0003,16'h004c,16'h001c,-16'h001b,16'h0027,-16'h0028,16'h0005,16'h002f,16'h001b,16'h0010,-16'h001e,-16'h0056,-16'h0049,16'h0034,16'h002b,16'h008a,-16'h006f,-16'h00ca,16'h0041,-16'h0033,-16'h0039,16'h0017,16'h0000,16'h0014,-16'h002a,16'h0025,-16'h0037,16'h002b,-16'h0016,16'h0027,16'h00ab,-16'h0086,16'h0025,-16'h00e8,-16'h001b,-16'h0010,16'h0000,-16'h005d,-16'h0034,-16'h0095,16'h003c,16'h0060,16'h0028,-16'h0089,16'h0004,-16'h010f,-16'h0014,16'h001c,-16'h0044,-16'h0079,16'h002c,16'h0070,16'h0058,-16'h0045,-16'h0061,16'h0010,16'h008c,16'h003a,16'h0045,16'h000b,-16'h001f,16'h0084,16'h0055,16'h0004,-16'h0018,-16'h0037,16'h0005,-16'h0057,16'h0012,-16'h0059,-16'h0073,16'h0028,16'h008f,-16'h0051,-16'h001c,-16'h0021,-16'h00c0,16'h0020,-16'h007f,16'h0029,-16'h0006,16'h0034,-16'h0062,-16'h0046,-16'h001d,-16'h0017,16'h0032,16'h0000,16'h0003,-16'h0090,16'h0026,16'h00aa,-16'h0003,16'h000a,16'h0023,16'h0053,-16'h0043,16'h000f,-16'h005e,16'h0042,16'h0004,-16'h001d,16'h000b,16'h0036,-16'h0009,-16'h009f,-16'h006d,16'h0032,-16'h0028,16'h003f,-16'h0006,16'h002a,16'h006a,16'h0033,16'h003f,-16'h0017,16'h0035,-16'h0015,-16'h007a,16'h008f,-16'h000a,16'h000e,16'h0042,16'h005f,16'h0047,-16'h0040,16'h0011,-16'h003d,16'h000e,16'h0035,-16'h001c,16'h0000,-16'h000d,-16'h009e,-16'h00a8,16'h0060,16'h001e,16'h002e,16'h003b,-16'h0036,16'h000a,-16'h0018,-16'h0025,16'h0037,-16'h000d,16'h0032,-16'h0041,-16'h002f,16'h000f,-16'h002e,16'h0030,-16'h0020,16'h0029,-16'h0079,16'h001a,16'h0098,-16'h0018,16'h004e,16'h001e,16'h0029,-16'h0093,-16'h0002,-16'h0059,16'h0038,-16'h0005,-16'h003e,-16'h004f,16'h0000,-16'h0002,-16'h0090,-16'h0060,16'h0018,-16'h002e,16'h0016,16'h003a,16'h001b,16'h006c,16'h0016,16'h0027,16'h0006,16'h0044,-16'h001c,-16'h0067,16'h00a4,-16'h001f,16'h002b,16'h002b,16'h001c,16'h002c,-16'h0015,16'h001c,-16'h0068,16'h0009,16'h0025,-16'h002a,16'h002c,-16'h002f,-16'h003d,-16'h00b9,16'h0063,16'h0000,16'h0041,16'h0004,-16'h000f,16'h002d,16'h001a,-16'h002c,16'h002c,16'h0014,-16'h0003,-16'h0056,-16'h001e,16'h001b,-16'h0018,16'h0035,-16'h001f,16'h0013,-16'h004d,-16'h003c,16'h007c,-16'h0046,16'h0056,16'h000a,16'h003f,-16'h009f,16'h0000,-16'h0089,16'h0035,16'h0044,-16'h0045,-16'h0046,16'h0007,16'h000c,-16'h00af,-16'h0040,16'h0039,16'h000c,-16'h001f,16'h0039,16'h0013,16'h0066,16'h0054,-16'h000a,16'h001c,16'h0005,-16'h0006,-16'h00a3,16'h0076,-16'h001a,16'h0030,16'h002e,16'h001d,16'h003a,16'h0016,-16'h0004,-16'h003d,-16'h0016,16'h0025,-16'h0027,16'h0027,16'h0009,-16'h0034,-16'h00e3,16'h004f,-16'h0003,16'h0026,16'h0004,-16'h0007,16'h003e,16'h003c,-16'h001b,16'h0037,16'h0001,16'h0010,-16'h0012,-16'h0058,16'h002e,-16'h0026,16'h0000,-16'h0020,16'h003b,-16'h0041,-16'h003e,16'h003e,-16'h002b,-16'h0011,-16'h0003,16'h0038,-16'h00ac,-16'h0003,-16'h00a7,16'h0000,16'h004a,-16'h0026,-16'h002d,16'h0003,-16'h0008,-16'h00c2,-16'h002f,16'h0015,16'h0001,-16'h0050,16'h0040,16'h001b,16'h003d,16'h0045,16'h0010,16'h0016,16'h0002,-16'h0038,-16'h00b2,16'h0094,16'h000e,16'h002c,16'h0028,16'h001c,16'h0050,16'h001a,-16'h0008,-16'h0058,16'h0003,16'h001d,-16'h000b,16'h0010,16'h000f,16'h0000,-16'h00dd,16'h0075,-16'h0016,16'h004a,-16'h0020,16'h0024,16'h0025,16'h0044,-16'h0021,16'h0032,16'h000d,16'h000d,-16'h0020,-16'h0059,16'h001f,-16'h0007,-16'h0002,-16'h0005,16'h0025,-16'h0013,-16'h0032,-16'h0011,-16'h0021,-16'h005c,16'h0020,-16'h0009,-16'h007b,16'h000a,-16'h00f5,-16'h0013,16'h0061,-16'h0062,-16'h005b,16'h0029,-16'h005d,-16'h0094,-16'h002e,16'h0025,16'h0018,-16'h0071,16'h002f,16'h000c,16'h0041,16'h0046,16'h002b,16'h0047,-16'h0023,-16'h0053,-16'h009c,16'h0079,-16'h0015,16'h0050,16'h0007,-16'h0014,16'h0088,16'h0056,-16'h001a,-16'h004e,16'h0022,16'h000e,-16'h003c,16'h0037,16'h0006,16'h0021,-16'h00c9,16'h0019,-16'h0021,16'h001b,16'h0009,16'h0025,16'h002b,16'h0048,16'h0027,16'h002f,16'h0046,-16'h0003,-16'h0008,-16'h009e,16'h0020,-16'h0030,-16'h0006,-16'h000b,16'h0024,-16'h004d,-16'h0021,-16'h0073,-16'h0001,-16'h00b3,16'h0051,16'h0004,-16'h0069,-16'h0029,-16'h00d9,-16'h001b,16'h002b,-16'h005a,-16'h0011,16'h0037,-16'h00b6,-16'h0058,16'h0000,16'h000f,16'h0023,-16'h007f,16'h001c,-16'h0036,16'h0041,16'h0011,16'h0054,16'h007c,-16'h0032,-16'h002d,-16'h007b,16'h0075,-16'h000d,16'h0055,-16'h0031,-16'h001d,16'h0087,16'h0045,-16'h0003,-16'h0045,16'h0033,16'h0011,-16'h001f,16'h001e,16'h0032,16'h0048,-16'h0075,-16'h0018,16'h0000,-16'h0002,16'h000e,16'h003c,16'h0029,16'h0060,16'h001d,16'h0025,16'h0003,16'h0008,16'h001f,-16'h0099,-16'h0004,-16'h0007,-16'h001c,-16'h0024,16'h0035,-16'h0048,-16'h0022,-16'h00b4,-16'h0004,-16'h0043,16'h0057,-16'h0015,-16'h0026,-16'h0033,-16'h00e7,-16'h0012,-16'h0016,-16'h0050,16'h0021,16'h005d,-16'h00b9,-16'h0076,-16'h0003,16'h0019,16'h0056,-16'h0045,16'h000d,-16'h0094,16'h003f,16'h000a,16'h009b,16'h0053,-16'h003b,-16'h001e,-16'h004e,16'h005f,-16'h004a,16'h0044,-16'h003f,-16'h001e,16'h0062,16'h000a,16'h0007,-16'h0051,16'h005a,16'h0005,-16'h0008,16'h002e,16'h0034,16'h0040,-16'h005c,-16'h0050,16'h0013,16'h0019,16'h0037,16'h002c,16'h001e,16'h006b,16'h0039,-16'h0003,-16'h0012,16'h0026,16'h0023,-16'h00a3,-16'h0009,-16'h000c,16'h0018,-16'h001f,16'h001e,-16'h0060,-16'h0046,-16'h00c2,-16'h0027,16'h004e,16'h0067,16'h000f,-16'h0001,-16'h002c,-16'h0088,-16'h000b,-16'h004d,-16'h0034,16'h0062,-16'h000f,-16'h0041,-16'h0061,16'h000f,16'h0020,16'h004e,-16'h0031,16'h002a,-16'h0083,16'h0043,-16'h0012,16'h00a3,16'h0016,-16'h002f,16'h0033,-16'h0031,16'h0033,-16'h004e,-16'h0002,-16'h0075,16'h0000,16'h004e,16'h0001,16'h002b,-16'h0065,16'h0051,-16'h0016,16'h000e,16'h003f,16'h000d,16'h0037,-16'h0074,-16'h0090,-16'h0010,16'h002c,16'h000d,16'h0031,16'h000c,16'h005b,16'h0019,-16'h0003,16'h0002,16'h0007,16'h0022,-16'h00b4,-16'h000b,16'h0036,16'h0001,-16'h0001,16'h001e,-16'h0056,-16'h001b,-16'h00f6,-16'h0030,16'h009b,16'h0047,16'h000a,16'h0029,-16'h004b,-16'h007b,-16'h001a,-16'h0076,16'h001f,16'h0035,-16'h0045,16'h0034,-16'h0048,-16'h0020,16'h0015,16'h0014,16'h0014,16'h001e,-16'h0063,16'h004f,-16'h0011,16'h0018,-16'h002c,-16'h0022,16'h0057,-16'h0021,16'h0036,-16'h0041,-16'h0045,-16'h00c5,16'h0004,16'h0060,-16'h0009,16'h0066,-16'h006f,16'h0007,-16'h0013,16'h0020,16'h0048,16'h001a,16'h0071,-16'h0055,-16'h00a7,16'h0002,16'h0008,16'h0008,16'h003f,16'h001a,16'h004c,16'h0021,16'h0000,16'h001a,16'h000c,16'h0031,-16'h0094,-16'h0005,16'h0019,16'h000b,16'h001c,16'h002e,-16'h0033,-16'h0016,-16'h0133,-16'h0024,16'h0048,16'h001a,16'h000b,16'h002f,-16'h0037,-16'h0051,-16'h0043,-16'h003a,16'h0069,16'h001a,-16'h0072,16'h0066,-16'h0046,-16'h0014,16'h0012,-16'h0018,16'h0025,16'h0017,16'h0019,16'h003b,16'h001e,-16'h0069,-16'h002a,-16'h001c,16'h0047,-16'h000f,16'h0038,16'h0016,-16'h0085,-16'h0114,16'h000c,16'h0077,-16'h0007,16'h002a,-16'h005a,16'h0017,-16'h0011,16'h003a,16'h003e,16'h005f,16'h0067,-16'h0058,16'h0009,16'h000a,-16'h000a,16'h0015,16'h0018,16'h000e,16'h0055,16'h0003,-16'h0029,16'h0009,-16'h0002,16'h001d,-16'h00a3,16'h002b,16'h0047,16'h0034,16'h002b,16'h0047,-16'h0029,16'h0000,-16'h0129,-16'h0022,-16'h0001,-16'h0028,16'h0012,16'h0029,-16'h0033,-16'h0026,-16'h0024,-16'h0009,16'h0061,16'h0015,-16'h0075,16'h0067,-16'h0044,-16'h001c,16'h0007,-16'h001e,16'h003b,16'h002b,16'h0083,16'h0047,16'h0051,-16'h008f,16'h004f,-16'h0002,16'h0008,-16'h000a,16'h0009,16'h002a,-16'h004c,-16'h012d,16'h003b,16'h0091,16'h001f,16'h0007,-16'h0079,16'h0031,-16'h001f,16'h0039,16'h003d,16'h0065,16'h005f,16'h0000,16'h0042,-16'h0024,16'h0013,16'h0039,-16'h001d,16'h0013,16'h005f,16'h0008,-16'h0016,16'h0011,-16'h0029,16'h003c,-16'h00a9,16'h003e,16'h002e,16'h0036,16'h0033,16'h0037,-16'h0001,16'h0030,-16'h00b6,16'h0005,-16'h0058,-16'h007d,-16'h0007,16'h001b,-16'h0032,-16'h0032,16'h0010,16'h0018,16'h0036,16'h0002,-16'h0077,16'h0042,-16'h002d,-16'h0008,16'h0019,-16'h0010,16'h0027,16'h0025,16'h007a,16'h0035,16'h003f,-16'h0046,16'h0056,16'h0013,-16'h005f,16'h0002,-16'h000e,16'h0050,-16'h0063,-16'h00ed,16'h0048,16'h0066,16'h0027,-16'h000c,-16'h005b,16'h000c,-16'h0028,16'h0040,16'h0022,16'h0050,16'h0059,16'h000e,16'h0075,-16'h0003,16'h0019,16'h0011,-16'h0010,16'h0011,16'h005a,16'h0005,-16'h0010,16'h0002,-16'h002c,16'h002b,-16'h00ac,16'h0056,16'h0025,16'h003a,16'h0003,16'h0021,-16'h0017,16'h0043,-16'h0020,16'h0012,-16'h0053,-16'h0064,-16'h000a,16'h003d,-16'h0012,-16'h001f,16'h0020,16'h000a,16'h0011,-16'h0004,-16'h0062,16'h0020,-16'h0035,-16'h001f,-16'h000f,16'h000a,-16'h0038,-16'h000d,16'h009c,16'h0043,16'h0048,16'h0037,16'h0024,16'h0009,-16'h0062,-16'h0003,-16'h0012,16'h0024,-16'h0057,-16'h0105,16'h0058,16'h0066,16'h0000,-16'h0019,-16'h003b,16'h0005,-16'h0009,16'h004e,16'h001e,16'h0020,16'h0039,16'h0043,16'h0048,16'h001d,16'h0011,16'h000c,-16'h0007,16'h0011,16'h0065,-16'h0001,16'h001a,16'h0001,-16'h0005,16'h0018,-16'h009e,16'h004a,16'h003e,16'h0051,-16'h001b,16'h0014,-16'h0004,16'h0040,16'h002f,16'h0013,-16'h002d,-16'h0065,16'h000b,16'h000a,-16'h000e,-16'h0035,16'h000b,16'h001b,16'h0028,-16'h002d,-16'h001e,-16'h004e,-16'h0065,16'h0033,-16'h0013,16'h003d,-16'h0051,-16'h0015,16'h0078,16'h0045,16'h0006,16'h005a,-16'h0063,16'h0002,16'h0006,16'h0009,-16'h0013,16'h003f,-16'h0053,-16'h009c,16'h006d,16'h001d,-16'h001c,-16'h0035,-16'h0054,16'h004d,-16'h000b,16'h002e,-16'h0007,16'h001d,16'h0036,16'h0070,16'h0030,16'h0011,16'h000f,16'h0026,-16'h0004,-16'h0026,16'h008a,16'h0022,-16'h0005,16'h0010,16'h002d,16'h000c,-16'h0094,16'h0060,16'h004c,16'h0030,-16'h0007,16'h0027,-16'h0019,16'h0019,16'h0036,16'h0032,16'h0002,-16'h000b,16'h000d,16'h0003,-16'h0014,-16'h0032,16'h0013,16'h0024,16'h000b,-16'h0015,-16'h0015,-16'h0077,-16'h005f,16'h003c,-16'h000f,16'h0060,-16'h0041,-16'h0027,16'h0075,16'h0053,-16'h003a,16'h0062,-16'h0086,-16'h001f,16'h000f,-16'h0003,-16'h0025,16'h0031,-16'h0036,-16'h001d,16'h0043,16'h0023,16'h003c,16'h0007,-16'h0046,16'h0031,16'h000c,16'h0018,-16'h001c,16'h0029,16'h0020,16'h007e,16'h000c,16'h0012,-16'h0001,16'h0010,16'h0016,-16'h0028,16'h00a0,16'h0034,16'h0010,16'h0003,-16'h0006,16'h0013,-16'h0080,16'h0072,16'h0039,16'h002e,16'h0002,16'h0027,-16'h003c,16'h0027,16'h004a,16'h0012,16'h003c,16'h0024,-16'h0003,16'h001a,-16'h0014,-16'h0031,16'h002f,-16'h000b,-16'h0007,-16'h001b,-16'h0019,-16'h0094,-16'h0039,16'h0033,-16'h000e,16'h002f,-16'h0046,-16'h002d,16'h006e,16'h0085,-16'h0071,16'h0057,-16'h004e,16'h0000,-16'h0004,16'h0008,-16'h000f,16'h0048,-16'h000d,16'h0028,16'h0012,16'h0040,16'h0022,-16'h001a,-16'h0026,16'h0016,16'h000e,16'h0010,-16'h0029,16'h0028,-16'h0027,16'h0079,-16'h001a,-16'h0018,-16'h0008,16'h0013,16'h002f,-16'h0026,16'h008c,16'h002c,16'h0020,16'h000f,-16'h0039,16'h000c,-16'h0076,16'h0035,16'h0042,16'h003b,-16'h0011,16'h003f,-16'h0012,16'h0013,16'h0031,16'h000e,16'h002b,16'h0044,-16'h0020,16'h0002,-16'h0021,-16'h0016,16'h0034,-16'h000e,16'h0012,-16'h001c,-16'h0016,-16'h002d,-16'h0030,16'h0031,-16'h0025,-16'h0005,-16'h0012,-16'h0026,16'h0033,16'h0072,-16'h00a4,16'h0057,16'h0011,-16'h0003,16'h0013,-16'h000c,-16'h000d,16'h002b,-16'h0010,16'h0070,16'h0007,16'h0023,16'h0015,16'h000a,16'h0000,-16'h000f,-16'h0008,-16'h0007,-16'h000e,16'h0026,-16'h003c,16'h0046,-16'h0043,16'h0002,16'h001f,16'h001d,16'h0045,-16'h0032,16'h0083,16'h0029,16'h002f,16'h0027,-16'h002b,16'h0018,-16'h0051,16'h0017,16'h003e,16'h0023,-16'h0025,16'h003a,-16'h0008,16'h0005,16'h0014,16'h0023,16'h0033,16'h0040,-16'h0026,16'h0000,-16'h004a,-16'h001d,16'h0006,-16'h0022,16'h000b,-16'h0002,16'h0007,-16'h0014,-16'h005f,16'h003f,-16'h001a,-16'h0010,16'h004f,16'h000b,-16'h0028,16'h0072,-16'h00af,16'h001d,16'h0042,16'h0008,-16'h0015,-16'h0007,-16'h0006,16'h000f,-16'h0020,16'h0075,-16'h0009,-16'h0006,16'h0012,16'h0011,-16'h001b,-16'h0010,-16'h0002,16'h0017,-16'h001f,16'h0015,-16'h0059,16'h0006,-16'h0021,16'h0015,16'h0020,16'h001b,16'h001d,-16'h003d,16'h007a,-16'h0004,16'h0011,16'h002c,-16'h0038,16'h002f,-16'h004e,-16'h0022,16'h0013,16'h0042,-16'h0041,16'h006e,16'h001f,-16'h000a,-16'h0033,16'h0004,16'h0032,16'h0043,-16'h0042,16'h000a,-16'h006b,-16'h0033,-16'h0014,16'h0002,16'h0016,16'h0018,-16'h001c,-16'h0024,-16'h0064,16'h001d,-16'h002d,-16'h0035,16'h0052,16'h001f,-16'h0046,16'h0054,16'h0008,16'h0014,16'h0057,-16'h0007,-16'h0001,16'h000d,16'h0013,-16'h0012,16'h0010,16'h0059,-16'h0014,-16'h0017,-16'h0013,-16'h0002,-16'h0007,-16'h0007,16'h000c,16'h003d,-16'h001e,16'h0000,-16'h003a,-16'h0003,16'h001f,16'h0039,16'h0002,16'h0028,16'h0000,-16'h003a,16'h0080,-16'h002e,16'h0018,-16'h000d,-16'h0046,16'h0022,-16'h0024,-16'h0039,16'h0016,16'h0058,-16'h0030,16'h0082,16'h0043,16'h0007,-16'h0009,-16'h000e,16'h0024,16'h0023,-16'h0028,16'h0021,-16'h0080,-16'h003d,-16'h0023,-16'h002a,16'h000f,16'h0005,-16'h0057,-16'h001b,-16'h0024,-16'h000e,-16'h002e,-16'h000c,16'h0050,16'h004a,-16'h0042,16'h003a,16'h0078,16'h0005,16'h002d,16'h000f,-16'h001c,16'h0016,16'h0031,-16'h0017,16'h0020,16'h003c,-16'h0004,-16'h001e,16'h000c,16'h0034,-16'h000a,-16'h0010,16'h000e,16'h003b,-16'h0020,16'h0003,-16'h002f,-16'h0023,16'h0024,16'h0055,16'h0005,16'h000e,16'h0005,-16'h0057,16'h0087,-16'h006e,16'h000c,16'h0012,-16'h0040,-16'h0001,-16'h0042,-16'h0097,16'h000c,16'h0028,-16'h002b,16'h004c,16'h0049,16'h002d,16'h0029,-16'h001a,-16'h000c,-16'h0033,-16'h001a,16'h0022,-16'h0087,-16'h0031,-16'h0021,-16'h0046,-16'h0004,-16'h0011,-16'h0056,16'h0040,16'h0010,-16'h0065,-16'h003a,16'h002e,16'h0063,16'h0044,-16'h000e,16'h001b,16'h008f,-16'h000c,-16'h0029,-16'h0014,-16'h005b,16'h0003,16'h0019,16'h0005,16'h003e,16'h003b,16'h000e,-16'h0018,16'h0020,16'h001e,16'h0025,-16'h002a,16'h0018,16'h001a,-16'h0009,16'h001f,-16'h0016,16'h0011,16'h0044,16'h0052,16'h000c,-16'h001b,-16'h000e,-16'h0011,16'h0071,-16'h0082,16'h001a,16'h002c,-16'h0079,-16'h0029,-16'h003b,-16'h00b2,16'h0008,16'h0023,-16'h003f,16'h0030,16'h0038,16'h0056,16'h0028,-16'h0016,-16'h001d,-16'h0064,-16'h0033,16'h0022,-16'h005c,-16'h004f,-16'h002a,-16'h00bd,-16'h0011,-16'h0018,-16'h0034,16'h005b,16'h000b,-16'h012d,-16'h0056,16'h000f,16'h0058,16'h0015,16'h000c,16'h0011,16'h0072,-16'h005c,-16'h0088,-16'h0026,-16'h005b,16'h0022,16'h0032,16'h001e,16'h0048,16'h0022,16'h0017,16'h0007,16'h003c,16'h0036,-16'h0009,16'h0004,16'h000d,16'h0005,-16'h001b,16'h0014,-16'h002b,16'h003d,16'h001d,16'h0020,16'h0020,-16'h0055,-16'h001c,16'h0018,16'h0040,-16'h008a,-16'h0017,16'h0023,-16'h0077,-16'h002b,-16'h0059,-16'h0079,16'h002e,16'h0024,-16'h0025,16'h002e,16'h004c,16'h0041,16'h0037,-16'h001a,-16'h001e,-16'h00a6,-16'h005a,16'h000b,-16'h0041,-16'h004b,-16'h0053,-16'h014c,-16'h0026,16'h002e,-16'h0034,16'h0024,16'h0002,-16'h01ed,-16'h0051,16'h0014,16'h0029,-16'h0057,16'h0049,16'h003d,16'h0025,-16'h0024,-16'h00c4,-16'h0031,16'h001d,16'h0024,16'h0014,16'h001e,16'h003c,16'h002b,16'h002c,16'h0000,16'h0043,16'h004f,16'h001c,-16'h0008,16'h004d,16'h000d,-16'h0009,16'h0020,-16'h0013,16'h0042,16'h0034,16'h0001,16'h0002,-16'h0046,-16'h0033,16'h0036,16'h007d,-16'h00c8,-16'h0023,16'h0018,-16'h0096,-16'h0014,-16'h004a,-16'h0054,-16'h000b,16'h0042,16'h0000,16'h0028,16'h000f,16'h0042,16'h002f,-16'h0002,16'h0000,-16'h00e1,-16'h0017,-16'h0042,-16'h006c,-16'h0026,-16'h003c,-16'h011f,-16'h003f,16'h0065,-16'h0025,16'h000c,-16'h0015,-16'h013d,-16'h0043,16'h0018,16'h0000,-16'h00a4,16'h0065,16'h002c,-16'h0079,-16'h000d,-16'h007a,-16'h003b,16'h0077,16'h004c,16'h0015,-16'h000a,16'h0036,16'h0018,16'h001a,16'h001a,16'h0022,16'h0046,-16'h0013,-16'h000e,16'h0036,16'h001c,16'h0005,-16'h000a,-16'h0003,16'h004d,16'h004c,16'h000a,16'h0019,-16'h002e,-16'h002b,16'h0056,16'h0062,-16'h0097,-16'h0019,16'h0015,-16'h008d,-16'h0004,-16'h003f,-16'h0033,-16'h0005,16'h000e,16'h0022,16'h002a,16'h0039,16'h0055,16'h0022,-16'h0027,-16'h0008,-16'h00d3,-16'h0019,-16'h002d,-16'h0053,-16'h000f,16'h0005,-16'h00ce,-16'h002e,16'h0059,-16'h003a,-16'h000c,-16'h0006,-16'h00c3,-16'h0033,-16'h0005,-16'h00bb,-16'h00be,16'h0085,16'h0030,-16'h0161,-16'h0016,16'h004b,-16'h0030,16'h008b,16'h000d,16'h001a,-16'h000c,16'h0051,16'h000e,-16'h0025,16'h0024,16'h0031,16'h0073,-16'h0011,-16'h0034,16'h0048,-16'h0007,16'h0013,16'h000e,16'h001d,16'h005a,16'h0030,16'h0020,16'h0021,-16'h0065,-16'h004f,16'h0050,16'h0067,-16'h0034,-16'h0008,16'h0003,-16'h0093,16'h0039,-16'h004a,-16'h000e,-16'h0014,16'h0011,16'h0041,-16'h0047,16'h0025,16'h005d,16'h0022,16'h0010,-16'h0001,-16'h0050,16'h0013,16'h0028,-16'h006a,-16'h0010,-16'h0008,-16'h0092,-16'h0010,16'h0030,-16'h0084,16'h000d,16'h0018,-16'h0096,-16'h0018,-16'h001e,-16'h0191,-16'h0078,16'h0072,16'h0031,-16'h0187,-16'h000e,16'h0070,-16'h000d,16'h003d,-16'h001f,16'h0044,16'h0022,16'h002f,16'h0048,16'h002d,16'h0045,16'h004e,16'h0051,16'h0002,-16'h002a,16'h006a,16'h0000,16'h002c,16'h0001,16'h0000,16'h000f,16'h003f,16'h0017,16'h002a,-16'h0017,-16'h0062,16'h0007,16'h006a,16'h0004,16'h0022,-16'h0013,-16'h0067,16'h0034,-16'h003e,-16'h001d,-16'h001f,-16'h0025,16'h0029,-16'h0071,16'h0028,16'h0049,16'h001e,16'h0029,16'h0010,16'h0032,-16'h0025,16'h0050,-16'h007b,16'h0002,-16'h003c,-16'h0049,-16'h0029,-16'h0020,-16'h00a1,16'h0001,16'h004d,-16'h005e,-16'h001b,-16'h004e,-16'h0156,-16'h002c,16'h0043,16'h0048,-16'h0112,-16'h0004,16'h0067,-16'h000d,-16'h0003,-16'h0030,16'h005d,16'h0016,16'h0024,16'h0066,16'h0035,16'h002b,16'h0034,16'h0051,16'h0004,-16'h000c,16'h0054,16'h0017,16'h0007,16'h000c,-16'h0033,-16'h0017,16'h0053,16'h0017,-16'h0001,-16'h0031,-16'h0050,-16'h0056,16'h007b,16'h0025,16'h0086,-16'h0037,-16'h00ac,16'h0029,-16'h0027,-16'h0027,-16'h0028,-16'h0029,-16'h000b,-16'h0064,16'h000e,-16'h001f,16'h004b,16'h000b,16'h003f,16'h007c,-16'h006f,16'h0036,-16'h00f1,-16'h0003,-16'h003c,-16'h0025,-16'h0072,-16'h003d,-16'h00a5,16'h0026,16'h005c,16'h002f,-16'h006a,-16'h0005,-16'h0131,-16'h0012,16'h0015,16'h0056,-16'h006e,16'h0021,16'h004c,16'h0014,-16'h003a,-16'h0067,16'h002c,16'h006e,16'h0029,16'h0032,16'h003f,-16'h0008,16'h0051,16'h0048,16'h0004,-16'h0033,-16'h0039,16'h001b,-16'h0066,-16'h0001,-16'h006a,-16'h0056,16'h0020,16'h009c,-16'h0059,-16'h0004,-16'h0025,-16'h00cf,16'h0045,-16'h006b,16'h0021,16'h0006,16'h0024,-16'h005d,-16'h0007,-16'h0035,-16'h002a,16'h003c,-16'h0008,16'h0017,-16'h00ab,16'h0027,16'h00ba,16'h001f,16'h0032,16'h0022,16'h0040,-16'h004f,-16'h000c,-16'h006a,16'h0050,-16'h0019,-16'h0007,16'h002e,16'h003b,16'h0021,-16'h00c6,-16'h0071,16'h0035,-16'h0038,16'h003c,16'h0015,16'h0056,16'h008a,16'h001e,16'h002e,-16'h000d,16'h0035,16'h0011,-16'h0080,16'h0075,-16'h0002,16'h002b,16'h000f,16'h0049,16'h0065,-16'h003c,16'h0015,-16'h0023,16'h001b,16'h0001,16'h0011,16'h0016,-16'h0026,-16'h0098,-16'h00ab,16'h0066,-16'h0021,16'h0012,16'h0035,-16'h004e,-16'h0049,16'h0000,-16'h0022,16'h0015,16'h0010,16'h0036,-16'h003a,16'h0001,-16'h0029,-16'h001d,16'h002c,16'h0009,16'h0010,-16'h00b3,-16'h0012,16'h00b6,16'h0000,16'h001f,16'h0022,16'h002d,-16'h00a6,16'h000d,-16'h006b,16'h0024,16'h002b,-16'h0046,-16'h002d,16'h0040,16'h000d,-16'h00f5,-16'h0059,16'h0016,-16'h0029,16'h0001,16'h0049,16'h0023,16'h0079,16'h0037,-16'h0002,16'h0008,16'h0028,-16'h0029,-16'h0082,16'h00a0,16'h000a,16'h0058,16'h000e,16'h0040,16'h004a,-16'h001e,16'h001e,-16'h002c,16'h0029,16'h0024,-16'h0026,16'h0012,-16'h0022,-16'h004b,-16'h00c7,16'h004a,-16'h0014,16'h000a,16'h002d,16'h0004,-16'h0033,16'h000b,-16'h0015,16'h0031,16'h0019,16'h0036,-16'h0017,16'h0026,16'h001c,-16'h0008,16'h0002,-16'h0015,16'h0021,-16'h00a2,-16'h0034,16'h0067,-16'h0001,-16'h0001,16'h0006,16'h003c,-16'h007d,16'h0024,-16'h00af,16'h001c,16'h0028,-16'h0034,-16'h004a,16'h001d,16'h0018,-16'h0123,-16'h0052,16'h0028,16'h000c,-16'h002c,16'h002b,16'h0028,16'h005e,16'h004b,-16'h0008,16'h0002,16'h0030,-16'h000d,-16'h0090,16'h009d,-16'h0008,16'h0054,16'h0002,16'h0003,16'h004e,-16'h000f,16'h0005,-16'h005f,16'h0026,16'h002a,-16'h0018,16'h001f,-16'h0021,-16'h0012,-16'h00eb,16'h005e,-16'h0023,16'h0031,-16'h0012,16'h0023,-16'h0021,16'h0007,-16'h0015,16'h001a,-16'h000d,16'h0043,16'h0010,16'h003f,16'h000e,-16'h0023,16'h001a,-16'h0015,16'h0028,-16'h0073,-16'h000d,-16'h0006,-16'h0033,-16'h0012,-16'h0008,16'h002c,-16'h0054,16'h0016,-16'h00cb,16'h0006,16'h0054,-16'h0045,-16'h0048,16'h0022,-16'h002a,-16'h012c,-16'h0072,16'h001b,16'h0002,-16'h0057,16'h0046,16'h0004,16'h0045,16'h0055,16'h0011,16'h0018,-16'h0004,-16'h002e,-16'h0084,16'h009c,-16'h0004,16'h003e,16'h001b,-16'h0006,16'h0077,16'h0000,-16'h000b,-16'h0093,16'h0029,16'h0017,-16'h0014,16'h0027,16'h0028,16'h0032,-16'h00f1,16'h0046,-16'h001b,16'h0034,16'h0003,16'h003a,-16'h001f,16'h0010,16'h001a,16'h000d,16'h0011,16'h0041,16'h0035,16'h0027,16'h002a,-16'h0033,-16'h0003,16'h000f,16'h001f,-16'h004c,16'h000d,-16'h0032,-16'h0023,-16'h0079,16'h0022,16'h0000,-16'h0039,16'h0015,-16'h012f,-16'h002c,16'h0067,-16'h0033,-16'h0043,16'h003d,-16'h00b6,-16'h00c2,16'h0000,16'h0020,16'h0003,-16'h008f,16'h0011,-16'h0014,16'h002f,16'h0043,16'h0056,16'h004b,-16'h000a,-16'h0045,-16'h0067,16'h00a9,16'h0001,16'h004f,16'h000e,-16'h000b,16'h0084,16'h001e,-16'h0033,-16'h00d0,16'h001e,16'h0011,-16'h000a,16'h002d,16'h0032,16'h0031,-16'h0097,16'h000c,-16'h0025,16'h0014,16'h000d,16'h0051,-16'h002a,16'h0030,16'h0035,16'h0011,16'h002a,16'h0020,16'h0003,16'h001c,16'h001d,-16'h0031,-16'h0007,16'h0022,16'h002d,-16'h0043,16'h000b,-16'h0043,-16'h0014,-16'h00c0,16'h003a,16'h000e,-16'h002a,16'h0006,-16'h0151,-16'h0029,16'h002a,-16'h0057,-16'h0011,16'h005c,-16'h00f1,-16'h0099,16'h0025,16'h002c,16'h0020,-16'h0071,16'h0019,-16'h005b,16'h0043,16'h0027,16'h0089,16'h0065,-16'h0029,-16'h0040,-16'h0049,16'h005b,-16'h000f,16'h003d,16'h0008,-16'h0003,16'h0080,16'h000c,16'h0005,-16'h0092,16'h0033,-16'h0008,16'h0010,16'h002b,16'h0020,16'h004e,-16'h0056,-16'h0025,-16'h002c,16'h0011,16'h0007,16'h004a,16'h0012,16'h0054,16'h0044,16'h0007,16'h0011,16'h0028,16'h000a,16'h001b,16'h0017,-16'h0036,-16'h000d,16'h001f,16'h0040,-16'h003e,16'h0021,-16'h009a,16'h0016,-16'h0040,16'h0070,-16'h0006,-16'h001f,-16'h000f,-16'h0153,16'h0000,-16'h001a,-16'h001f,16'h0020,16'h0068,-16'h0066,-16'h0087,16'h001e,16'h0046,16'h005c,-16'h0022,16'h0001,-16'h00b2,16'h005e,-16'h0026,16'h009c,16'h0052,16'h0000,-16'h0031,-16'h0036,16'h003b,-16'h0034,-16'h0003,16'h0025,16'h0001,16'h004f,-16'h0003,16'h0020,-16'h007b,16'h003e,-16'h0016,16'h0028,16'h002f,16'h0004,16'h0045,-16'h0028,-16'h002f,-16'h000f,16'h0023,16'h0013,16'h0058,16'h0005,16'h0050,16'h004a,-16'h0037,-16'h0007,16'h0030,16'h0025,-16'h000c,-16'h0006,-16'h001d,-16'h0004,16'h0009,16'h002e,-16'h0024,16'h0029,-16'h00df,16'h0012,16'h001b,16'h003d,16'h000a,-16'h000e,-16'h0026,-16'h015a,16'h001a,-16'h005e,16'h0001,16'h0043,16'h0037,16'h000f,-16'h0072,16'h0040,16'h0053,16'h005c,16'h0028,16'h0028,-16'h00a0,16'h0040,-16'h0022,16'h0077,-16'h000d,-16'h000f,16'h003d,-16'h0021,16'h001e,-16'h0060,-16'h003a,16'h0030,16'h0006,16'h005a,-16'h0009,16'h005e,-16'h0077,16'h0045,-16'h0033,16'h0022,16'h0001,16'h0002,16'h0085,-16'h0026,-16'h0084,-16'h0007,16'h001a,16'h002a,16'h001c,16'h000b,16'h0047,16'h001c,-16'h0037,16'h0004,-16'h0005,16'h0046,16'h0005,-16'h0019,-16'h0016,-16'h0003,-16'h000d,16'h004f,-16'h0019,16'h003e,-16'h013d,16'h0013,16'h005d,16'h0000,16'h0002,16'h0006,-16'h0027,-16'h0183,-16'h002e,-16'h0076,16'h0065,16'h0029,-16'h001f,16'h0058,-16'h0083,16'h0029,16'h005d,16'h0038,16'h003e,16'h001b,-16'h004c,16'h006e,-16'h0001,-16'h002e,-16'h004f,-16'h000f,16'h0097,16'h0002,-16'h000e,-16'h0045,-16'h00af,-16'h0019,16'h0020,16'h0074,16'h0007,16'h0058,-16'h0074,16'h0010,16'h000a,16'h003f,16'h0025,16'h0038,16'h0089,-16'h003d,-16'h008c,16'h0006,16'h0021,16'h0008,16'h000f,16'h0021,16'h0044,16'h004b,-16'h001f,16'h001a,16'h000c,16'h004a,-16'h001c,-16'h0003,16'h000c,-16'h0002,16'h001f,16'h0032,16'h0010,16'h0033,-16'h014c,16'h0003,16'h0040,-16'h0011,16'h0008,16'h0028,-16'h0038,-16'h0137,-16'h0034,-16'h001b,16'h0083,16'h001a,-16'h006a,16'h0062,-16'h009a,16'h0007,16'h0057,-16'h001d,16'h0050,16'h0013,16'h0028,16'h006e,16'h004a,-16'h005c,16'h001b,-16'h002a,16'h004b,-16'h0005,-16'h002e,16'h002a,-16'h005e,-16'h0075,16'h0041,16'h0096,16'h0002,16'h0041,-16'h0054,16'h0015,-16'h0011,16'h0038,16'h0006,16'h0075,16'h008c,16'h0017,-16'h0032,16'h0013,16'h0010,16'h0015,16'h0019,16'h000d,16'h0043,16'h003a,-16'h0042,16'h0011,-16'h0004,16'h001b,-16'h002a,16'h000d,16'h001a,-16'h000e,16'h001d,16'h004b,16'h0047,16'h0057,-16'h00d7,16'h0023,-16'h000d,-16'h0043,16'h0007,16'h0041,-16'h0060,-16'h00db,-16'h0028,16'h001e,16'h0071,-16'h000c,-16'h0064,16'h005a,-16'h0058,-16'h001a,16'h0050,-16'h0027,16'h005b,16'h0030,16'h007e,16'h0058,16'h0078,-16'h008f,16'h0048,-16'h0019,-16'h0032,16'h0020,-16'h0045,16'h003b,16'h0001,-16'h00a1,16'h005c,16'h0091,16'h0000,16'h002e,-16'h0061,16'h0028,-16'h0008,16'h0036,16'h0012,16'h0061,16'h0054,16'h0040,16'h0031,-16'h000f,16'h002a,-16'h0007,16'h0009,-16'h001a,16'h004f,16'h002b,-16'h002a,16'h0005,-16'h0001,16'h0014,-16'h003f,16'h0010,16'h0012,-16'h000e,16'h003a,16'h003a,16'h004e,16'h0060,-16'h0019,16'h0038,-16'h006f,-16'h004e,16'h0005,16'h001c,-16'h004d,-16'h00c7,16'h0002,16'h002c,-16'h0017,16'h000b,-16'h0072,16'h0036,-16'h0076,-16'h001e,16'h0056,-16'h000d,16'h0024,16'h0023,16'h0089,16'h005a,16'h002d,-16'h003d,16'h003c,16'h000a,-16'h006b,16'h0024,-16'h003f,16'h0029,16'h0003,-16'h00c5,16'h0032,16'h0065,-16'h000e,16'h000b,-16'h006b,16'h003b,-16'h0015,16'h0019,16'h0003,16'h0064,16'h0056,16'h0061,16'h0059,-16'h001c,16'h0032,16'h0010,-16'h0008,-16'h0025,16'h004f,16'h001b,-16'h001d,-16'h0008,16'h0027,16'h0024,-16'h0053,16'h0019,16'h0008,16'h0018,16'h000e,16'h0005,16'h0017,16'h004b,16'h0061,16'h001d,-16'h0047,-16'h005f,-16'h0005,16'h0025,-16'h004f,-16'h0099,16'h000a,16'h0017,-16'h0008,16'h0002,-16'h0064,-16'h0009,-16'h0080,-16'h0016,16'h0065,16'h0037,-16'h0034,16'h0000,16'h009d,16'h0077,16'h0040,16'h003e,-16'h0018,16'h000a,-16'h009f,16'h0024,-16'h0047,16'h0035,-16'h000b,-16'h0100,16'h0047,16'h0063,-16'h002f,-16'h0011,-16'h004e,16'h0035,-16'h0009,16'h0018,16'h0013,16'h003b,16'h0017,16'h0075,16'h004f,16'h0008,16'h0027,-16'h0001,-16'h0026,-16'h002f,16'h003c,16'h0002,-16'h0009,-16'h0008,16'h002d,16'h002d,-16'h0052,16'h003f,16'h000b,16'h0027,-16'h0010,16'h0023,16'h004c,16'h000f,16'h0082,16'h0034,-16'h003a,-16'h006f,-16'h0016,16'h000d,-16'h0059,-16'h0089,-16'h000d,16'h0001,16'h002c,-16'h001d,-16'h0044,-16'h008d,-16'h007a,16'h0026,16'h0065,16'h0038,-16'h0059,16'h0011,16'h0056,16'h0094,16'h002f,16'h005c,-16'h0051,16'h0009,16'h0000,16'h0007,-16'h0052,16'h0022,-16'h0033,-16'h00bf,16'h004e,16'h0027,-16'h001a,-16'h002b,-16'h004c,16'h0042,16'h0003,16'h0008,-16'h0016,16'h000d,-16'h001e,16'h008a,16'h004a,16'h000f,16'h002b,16'h001b,-16'h0025,-16'h0045,16'h002e,-16'h0038,-16'h0009,-16'h000d,16'h004b,16'h0007,-16'h0051,16'h0042,16'h0019,16'h0025,16'h000f,16'h0019,16'h0015,-16'h0006,16'h0088,16'h003e,-16'h0011,-16'h0033,-16'h000a,-16'h0021,-16'h006d,-16'h007a,-16'h0010,16'h0036,16'h001c,-16'h0019,-16'h0017,-16'h0089,-16'h0076,16'h002a,16'h0061,16'h0054,-16'h0050,-16'h0016,16'h0046,16'h0087,-16'h0023,16'h0045,-16'h0069,-16'h0002,16'h0012,16'h0012,-16'h005a,16'h001a,16'h0004,-16'h0098,16'h0032,16'h0046,16'h0003,16'h0010,-16'h0035,16'h003b,-16'h0008,-16'h0012,-16'h0004,16'h0040,-16'h0029,16'h0079,16'h000d,16'h0003,-16'h0002,16'h0011,16'h001d,-16'h0024,16'h0047,-16'h0012,16'h0002,-16'h0022,16'h0063,16'h002a,-16'h0045,16'h0033,-16'h0021,16'h0012,16'h0025,16'h0026,16'h0028,16'h0004,16'h0089,16'h0021,16'h0004,16'h0021,-16'h0004,16'h0004,-16'h0066,-16'h007b,16'h0016,16'h0016,16'h0009,-16'h0012,16'h0006,-16'h0084,-16'h0050,16'h004b,16'h007b,16'h001d,-16'h0074,-16'h0046,16'h002e,16'h0090,-16'h0077,16'h005b,-16'h0047,-16'h0007,16'h001c,-16'h0009,-16'h0041,16'h0030,16'h000d,-16'h004b,16'h0005,16'h004a,-16'h0006,-16'h001b,-16'h0012,16'h0036,-16'h001f,-16'h001b,16'h0007,16'h0040,-16'h0040,16'h0073,-16'h0034,-16'h000b,-16'h000b,16'h0005,16'h0012,-16'h0021,16'h005e,-16'h001e,16'h000f,-16'h0018,16'h0022,16'h0022,-16'h0049,16'h004c,-16'h0004,16'h001b,16'h0018,16'h0026,-16'h001c,16'h000e,16'h0049,16'h0032,16'h0022,16'h0026,16'h000e,-16'h0003,-16'h0076,-16'h0064,16'h0011,16'h0007,-16'h0019,-16'h0029,-16'h0004,-16'h0035,-16'h005d,16'h0043,16'h0075,16'h0002,-16'h0037,-16'h002e,-16'h0057,16'h0074,-16'h00ad,16'h004a,16'h0007,-16'h0018,-16'h0002,16'h0001,-16'h003c,16'h000a,16'h0011,16'h0019,-16'h0003,16'h0042,-16'h000c,16'h0004,-16'h000a,16'h0031,-16'h0002,16'h0002,-16'h0015,16'h001c,-16'h0052,16'h0037,-16'h009a,16'h0006,16'h0019,16'h0001,16'h002d,-16'h0042,16'h0050,16'h0009,16'h0029,-16'h000c,16'h003a,16'h0010,-16'h0038,16'h0053,16'h001b,16'h0034,-16'h0008,16'h001d,16'h0011,-16'h0028,16'h0010,16'h004b,16'h002c,16'h001c,-16'h0014,16'h0013,-16'h0074,-16'h005d,16'h000a,-16'h001d,-16'h0008,16'h0012,16'h0004,-16'h000d,-16'h004b,16'h0051,16'h0065,-16'h0007,16'h0037,16'h0016,-16'h0083,16'h0073,-16'h0089,16'h0015,16'h001a,-16'h0023,-16'h0003,16'h0004,16'h0007,16'h001a,16'h0000,16'h0056,-16'h001d,-16'h0001,-16'h0008,16'h0000,16'h0015,16'h001a,-16'h000a,16'h001c,16'h0001,16'h0002,-16'h0044,-16'h0014,-16'h0064,16'h001c,16'h0012,16'h0001,16'h001f,-16'h0044,16'h005a,-16'h0030,16'h0034,-16'h000b,16'h001b,16'h0016,-16'h0025,16'h0035,16'h001f,16'h005b,-16'h0025,16'h0075,16'h000a,-16'h0044,-16'h0020,16'h0029,16'h002b,16'h000b,16'h0003,16'h0030,-16'h0069,-16'h0084,16'h000c,-16'h001d,16'h0004,16'h0010,-16'h0013,16'h0003,-16'h0067,16'h0034,16'h0039,-16'h002e,16'h0059,16'h0017,-16'h006b,16'h005f,16'h003c,16'h000a,16'h003d,-16'h0003,-16'h0003,16'h0016,16'h0042,-16'h0016,16'h0026,16'h0052,-16'h000c,-16'h001d,-16'h0020,-16'h0025,16'h0005,16'h000f,-16'h0030,16'h003a,-16'h000e,-16'h000b,-16'h002d,-16'h002e,-16'h002e,16'h0024,16'h000a,16'h0011,16'h0039,-16'h0034,16'h0071,-16'h0045,16'h001d,-16'h0009,16'h0015,16'h0024,-16'h0006,16'h001b,16'h0035,16'h003e,-16'h003f,16'h006a,16'h000a,-16'h000a,-16'h0023,16'h000f,16'h0024,16'h0000,-16'h0018,16'h004b,-16'h0074,-16'h005c,-16'h0034,-16'h0041,16'h0000,16'h001b,-16'h0029,16'h002b,-16'h0034,-16'h0010,16'h0042,-16'h0011,16'h0061,16'h002c,-16'h0063,16'h0065,16'h005b,16'h0025,16'h0016,-16'h0013,-16'h0019,16'h0023,16'h0045,-16'h0011,16'h0009,16'h0059,-16'h0009,-16'h000f,16'h0003,-16'h000c,16'h000a,-16'h0016,-16'h0006,16'h0061,16'h0004,-16'h0012,-16'h0022,-16'h003f,-16'h0015,16'h0065,16'h000e,-16'h000d,16'h0016,-16'h0016,16'h0060,-16'h004d,16'h0014,-16'h000b,-16'h0015,16'h0002,-16'h0014,-16'h0041,16'h001d,16'h0015,-16'h0030,16'h0052,16'h000d,16'h0015,-16'h0018,16'h001d,-16'h0004,-16'h0030,-16'h0016,16'h0023,-16'h0089,-16'h0072,-16'h0043,-16'h004c,-16'h0015,16'h0006,-16'h003c,16'h0049,-16'h000c,-16'h0070,-16'h0002,16'h0014,16'h0072,16'h002e,-16'h0038,16'h0058,16'h007a,-16'h002c,-16'h0042,-16'h000e,-16'h0043,16'h001b,16'h0041,16'h0003,16'h004e,16'h0068,16'h0012,16'h001c,-16'h0006,16'h0019,16'h001a,-16'h002c,16'h0015,16'h0010,16'h0012,-16'h000d,-16'h0028,-16'h0009,-16'h000f,16'h0039,16'h0019,-16'h004b,16'h0013,16'h0008,16'h0040,-16'h005f,16'h000d,16'h000a,-16'h0006,-16'h000c,16'h000c,-16'h007b,16'h0037,16'h0003,-16'h000d,16'h0034,16'h0023,16'h0049,-16'h0001,16'h001c,-16'h0023,-16'h0046,-16'h0016,16'h0009,-16'h006a,-16'h005c,-16'h0040,-16'h0064,16'h0008,-16'h0006,-16'h0025,16'h0070,-16'h000b,-16'h01b3,-16'h0010,16'h0015,16'h0059,16'h0027,16'h0010,16'h005e,16'h008d,-16'h007e,-16'h0080,-16'h0037,-16'h0028,16'h0011,16'h0020,16'h0025,16'h003e,16'h0044,16'h003c,16'h0011,16'h0001,16'h002f,16'h0022,16'h000a,16'h002f,16'h0022,-16'h000e,16'h001b,-16'h0001,16'h0016,-16'h001a,16'h0029,16'h0015,-16'h0058,16'h0015,16'h0010,16'h0054,-16'h0064,-16'h0013,16'h000b,-16'h001b,-16'h0019,-16'h000c,-16'h008e,16'h001e,16'h000f,16'h0000,16'h0028,16'h0009,16'h006b,16'h0015,-16'h0003,16'h0003,-16'h0072,-16'h0025,-16'h0004,-16'h008f,-16'h005d,-16'h004c,-16'h010f,-16'h0002,16'h0034,-16'h001e,16'h0035,-16'h0023,-16'h025f,-16'h0026,16'h0021,16'h002e,-16'h0035,16'h0046,16'h004a,16'h000d,-16'h002b,-16'h004a,-16'h0031,16'h001d,16'h0027,16'h0023,-16'h002e,16'h0033,16'h002c,16'h003d,16'h0024,-16'h0011,16'h004d,16'h001d,16'h001c,16'h002f,16'h0016,-16'h000d,16'h0002,16'h0012,16'h002f,16'h001f,16'h0020,-16'h0008,-16'h0068,-16'h002d,16'h004a,16'h0064,-16'h0070,-16'h0021,16'h000b,-16'h0058,-16'h0012,-16'h0012,-16'h00a6,-16'h0009,16'h0015,16'h002f,16'h0007,16'h0007,16'h0065,16'h004e,16'h0002,-16'h0003,-16'h00c2,-16'h0015,-16'h0023,-16'h0088,-16'h0054,-16'h0024,-16'h012f,16'h000f,16'h0059,-16'h000c,16'h000e,-16'h004d,-16'h0130,-16'h0013,16'h0022,16'h0013,-16'h00af,16'h004f,16'h0050,-16'h00a2,16'h0008,-16'h0008,-16'h0046,16'h0071,16'h003d,16'h0010,-16'h0019,16'h0029,16'h002a,16'h003e,16'h0027,16'h001d,16'h0057,16'h000f,16'h001e,16'h0053,16'h0009,-16'h0011,-16'h000d,16'h0016,16'h0042,16'h004f,16'h0011,16'h0029,-16'h0036,-16'h007d,16'h006b,16'h0071,-16'h009b,-16'h0006,-16'h0012,-16'h0066,-16'h0017,16'h0003,-16'h005a,-16'h002f,16'h001b,16'h0019,-16'h0028,16'h005a,16'h0063,16'h0046,-16'h0001,-16'h0012,-16'h00be,-16'h0008,-16'h0021,-16'h0075,-16'h0053,-16'h0001,-16'h00fe,-16'h0007,16'h0063,-16'h004b,-16'h001d,-16'h0043,-16'h00bb,-16'h0036,-16'h0034,-16'h00e0,-16'h0093,16'h0074,16'h0041,-16'h0172,16'h0003,16'h0034,-16'h0041,16'h0069,16'h000d,16'h001a,-16'h0001,16'h0027,16'h001d,16'h001c,16'h0048,16'h003c,16'h0061,-16'h0022,-16'h0006,16'h003f,16'h0000,-16'h001d,16'h0008,16'h000d,16'h002d,16'h0038,16'h004b,16'h0045,-16'h0049,-16'h008b,16'h0057,16'h005b,-16'h007b,-16'h000e,-16'h0006,-16'h0045,16'h0019,-16'h0022,-16'h002d,-16'h0046,-16'h001f,16'h0041,-16'h006c,16'h0047,16'h0047,16'h004c,16'h001f,-16'h0005,-16'h004e,16'h0001,16'h0025,-16'h007d,-16'h0030,16'h0003,-16'h0089,-16'h0028,-16'h001c,-16'h008b,-16'h000d,-16'h0020,-16'h00af,-16'h001b,-16'h004d,-16'h01da,-16'h0056,16'h0048,16'h0053,-16'h0158,16'h0017,16'h0068,-16'h001c,16'h001a,-16'h0016,16'h0053,-16'h0014,16'h0016,16'h0044,16'h004a,16'h0068,16'h0017,16'h003f,-16'h0018,16'h0003,16'h003d,16'h0006,16'h000c,16'h0004,16'h001a,16'h0005,16'h0059,16'h001d,16'h0026,-16'h0037,-16'h005c,-16'h0013,16'h0067,-16'h002b,16'h0032,-16'h0002,-16'h003b,16'h0026,-16'h0032,-16'h001e,-16'h0063,-16'h0020,-16'h0011,-16'h009a,16'h001a,16'h0054,16'h0051,16'h0030,16'h0025,16'h001a,-16'h0012,16'h001a,-16'h009f,-16'h0022,-16'h0049,-16'h0053,-16'h0041,-16'h0043,-16'h00b6,-16'h000f,16'h0001,-16'h0029,-16'h001c,-16'h0044,-16'h0189,-16'h0041,16'h0014,16'h0069,-16'h0112,16'h0046,16'h0062,-16'h0027,-16'h000d,-16'h000c,16'h0061,-16'h001a,16'h0014,16'h0047,16'h0068,16'h0043,16'h0010,16'h0033,-16'h000e,16'h000f,16'h0045,16'h002e,-16'h0006,-16'h0009,-16'h001c,-16'h0025,16'h0051,16'h0028,-16'h0018,-16'h0013,-16'h003a,-16'h005f,16'h0079,16'h000c,16'h005d,-16'h0021,-16'h006f,16'h001c,-16'h0016,-16'h004a,-16'h0034,-16'h002a,-16'h0043,-16'h0096,16'h0010,-16'h001e,16'h0057,16'h0042,16'h0057,16'h0040,-16'h0043,-16'h0006,-16'h0107,-16'h0002,-16'h002e,-16'h0030,-16'h0081,-16'h004a,-16'h00bb,-16'h0003,16'h0025,16'h003b,-16'h0048,-16'h000d,-16'h0123,-16'h001f,16'h0010,16'h0075,-16'h0070,16'h001e,16'h0049,16'h000d,-16'h0028,-16'h0038,16'h003c,16'h0025,16'h001b,16'h000c,16'h007f,-16'h0018,-16'h0001,16'h0005,-16'h0019,-16'h0024,-16'h0018,16'h001d,-16'h0028,16'h0003,-16'h0042,-16'h0052,16'h001f,16'h008a,-16'h0076,-16'h0034,-16'h0016,-16'h00f3,16'h0079,-16'h0088,16'h0032,-16'h0012,16'h0034,-16'h001c,-16'h0009,-16'h000d,-16'h0018,16'h0033,16'h0000,16'h0017,-16'h008e,16'h0031,16'h0090,16'h004e,16'h003d,16'h0016,16'h0045,-16'h0042,16'h0006,-16'h0058,16'h002c,-16'h0013,-16'h0027,16'h005b,16'h003c,16'h0021,-16'h00c6,-16'h0061,16'h0001,-16'h004d,16'h0037,16'h005a,16'h0030,16'h0082,16'h0002,16'h0000,-16'h0021,16'h0012,-16'h0011,-16'h0046,16'h0085,16'h000f,16'h0014,16'h004e,16'h003a,16'h0061,-16'h002e,16'h0006,-16'h000f,16'h004e,-16'h0045,16'h0018,16'h000e,-16'h004a,-16'h0059,-16'h00c7,16'h002f,-16'h002c,16'h0016,16'h0034,-16'h0033,-16'h00a0,-16'h0037,-16'h003f,16'h0010,16'h0014,16'h003c,16'h0018,16'h003d,-16'h001c,-16'h0011,16'h002d,-16'h000e,16'h0020,-16'h009a,-16'h0015,16'h0085,16'h0021,16'h002d,16'h0004,16'h003f,-16'h0046,16'h0033,-16'h0041,16'h0011,16'h0017,-16'h0043,-16'h001f,16'h0024,-16'h0016,-16'h0126,-16'h0079,16'h0012,-16'h0052,16'h001b,16'h004b,16'h0045,16'h0075,16'h004f,16'h0007,16'h000f,16'h0031,-16'h001f,-16'h0038,16'h00bc,16'h0019,16'h0033,16'h0036,16'h0053,16'h0050,-16'h0022,16'h001c,-16'h000b,16'h004f,-16'h0017,-16'h0023,16'h002d,-16'h0037,-16'h003d,-16'h00ce,16'h0035,-16'h003b,16'h0006,16'h001a,-16'h001b,-16'h00d4,-16'h001d,-16'h000b,16'h0006,16'h0000,16'h0056,16'h0022,16'h005f,16'h001b,-16'h002a,16'h0000,-16'h0014,16'h0023,-16'h00c1,-16'h001b,16'h002c,16'h0029,-16'h001a,-16'h000a,16'h001c,-16'h0017,16'h003c,-16'h005e,-16'h0007,16'h0038,-16'h006d,-16'h002f,16'h0010,-16'h0048,-16'h014f,-16'h0074,16'h0011,-16'h0055,16'h0007,16'h005b,16'h0010,16'h004c,16'h004e,16'h0011,16'h0000,16'h0034,-16'h0006,-16'h004e,16'h00b0,16'h002a,16'h002d,16'h000f,16'h0038,16'h005e,-16'h0016,16'h0014,-16'h005d,16'h0028,16'h0016,-16'h002f,16'h0011,-16'h0010,16'h0014,-16'h00d3,16'h004e,-16'h0031,16'h000f,16'h0015,16'h0000,-16'h00cb,-16'h0020,16'h0024,16'h0023,-16'h001a,16'h006d,16'h0049,16'h0096,16'h0016,-16'h0025,16'h0020,16'h002d,16'h001a,-16'h0085,16'h0004,-16'h006e,16'h001d,-16'h003b,16'h0000,-16'h0012,16'h000b,16'h001d,-16'h007b,-16'h0036,16'h0066,-16'h0062,-16'h003d,16'h0022,-16'h008c,-16'h0189,-16'h0059,16'h0005,-16'h002c,-16'h0036,16'h005f,16'h0007,16'h0014,16'h0034,16'h0039,16'h002b,16'h001c,16'h0006,-16'h0039,16'h009a,-16'h0009,16'h000f,16'h000c,-16'h0003,16'h007d,-16'h0013,-16'h0014,-16'h007b,16'h0038,16'h002a,-16'h0008,16'h002e,-16'h0006,16'h0033,-16'h00d9,16'h0056,-16'h0022,16'h0026,16'h0006,16'h0065,-16'h00f0,16'h0011,16'h0044,16'h001a,16'h000b,16'h0065,16'h002a,16'h009a,16'h000f,-16'h0023,-16'h0008,16'h0032,16'h002e,-16'h0046,16'h0022,-16'h0092,16'h000c,-16'h0073,16'h001b,16'h0011,16'h0017,16'h0020,-16'h00bd,-16'h0041,16'h005b,-16'h0048,-16'h0035,16'h0058,-16'h00c7,-16'h00fa,-16'h0022,16'h0027,16'h0007,-16'h0057,16'h002f,-16'h0023,16'h000b,16'h0027,16'h005e,16'h0036,-16'h0003,-16'h002c,-16'h003d,16'h006c,16'h000c,16'h000d,16'h000a,-16'h0003,16'h008b,-16'h0011,-16'h000d,-16'h00a9,16'h003e,16'h0017,16'h0029,16'h0028,16'h0001,16'h0026,-16'h006d,16'h0000,-16'h002c,16'h0000,-16'h0001,16'h007e,-16'h00e4,16'h0026,16'h003d,16'h0026,16'h0023,16'h0043,16'h0010,16'h0084,16'h0033,-16'h0040,-16'h0008,16'h0033,16'h001f,-16'h0056,16'h004d,-16'h00b0,16'h004a,-16'h00a1,16'h005c,16'h0001,16'h0011,16'h0020,-16'h00d9,-16'h0004,16'h001f,-16'h0064,16'h0004,16'h007f,-16'h00be,-16'h00b1,16'h000d,16'h0022,16'h0048,-16'h003f,16'h0023,-16'h00b5,16'h0008,-16'h0005,16'h008b,16'h005d,-16'h0004,-16'h001b,-16'h0022,16'h0047,-16'h002e,16'h001b,16'h000a,16'h0018,16'h007a,-16'h0009,-16'h0021,-16'h00a7,16'h0002,-16'h000c,16'h0034,16'h0023,-16'h0013,16'h0044,-16'h003d,-16'h001b,-16'h001f,-16'h001a,-16'h0016,16'h0089,-16'h0084,16'h0044,16'h004e,16'h0007,16'h001d,16'h0034,16'h0002,16'h0097,16'h0045,-16'h0054,16'h000a,16'h003a,16'h0017,-16'h0022,16'h0045,-16'h00aa,16'h003c,-16'h0057,16'h005c,-16'h000e,-16'h0028,16'h0020,-16'h00e6,16'h0001,-16'h0019,-16'h0021,16'h003f,16'h007f,-16'h0015,-16'h008b,16'h003f,16'h002d,16'h005b,16'h0007,16'h0018,-16'h00dc,16'h001f,-16'h004b,16'h00a7,16'h0027,-16'h001c,16'h0017,16'h0002,16'h003e,-16'h004e,-16'h0019,16'h002d,16'h002a,16'h003b,-16'h000f,16'h0022,-16'h0089,16'h0024,-16'h0004,16'h0027,16'h0014,-16'h0009,16'h0050,-16'h0006,-16'h0049,-16'h0022,-16'h0009,-16'h000a,16'h0083,-16'h006f,16'h0055,16'h0040,-16'h0020,16'h000b,16'h000e,-16'h0007,16'h00a2,16'h0028,-16'h004e,-16'h0013,16'h0016,16'h000d,-16'h000d,16'h0075,-16'h00bc,16'h004d,16'h002e,16'h002b,-16'h000b,16'h000c,16'h0027,-16'h00ec,-16'h000f,-16'h0046,16'h002c,16'h0024,16'h0060,16'h0064,-16'h007c,16'h0036,16'h002a,16'h0058,16'h0020,16'h0020,-16'h00a2,16'h0023,-16'h002f,16'h0055,-16'h003d,-16'h0003,16'h006c,-16'h0002,-16'h000f,-16'h0059,-16'h0043,16'h006b,16'h002b,16'h0032,16'h0024,16'h0063,-16'h007c,16'h0002,-16'h0024,16'h0043,16'h0011,16'h0000,16'h006e,16'h000b,-16'h007d,16'h002d,16'h0020,16'h001b,16'h0049,-16'h0035,16'h0039,16'h0042,-16'h0018,-16'h0002,16'h000e,16'h000e,16'h0095,16'h0010,-16'h0023,16'h0000,16'h000f,16'h0027,16'h0012,16'h0095,-16'h00eb,16'h0057,16'h0048,-16'h0004,16'h000c,16'h0001,16'h0019,-16'h0118,-16'h0004,-16'h0061,16'h0053,16'h0029,16'h001a,16'h006f,-16'h0089,16'h0028,16'h0052,16'h000b,16'h0049,16'h0005,-16'h0025,16'h0035,16'h002d,-16'h000c,-16'h0056,-16'h0016,16'h0099,-16'h0011,-16'h0033,-16'h004c,-16'h0094,16'h0054,16'h0021,16'h006f,16'h002f,16'h006c,-16'h0096,16'h0012,-16'h0018,16'h0051,16'h0006,16'h0041,16'h0089,16'h0033,-16'h0069,16'h003b,16'h003b,16'h0021,16'h0045,-16'h0038,16'h0030,16'h007b,-16'h0033,16'h0021,-16'h0005,16'h0026,16'h00a1,-16'h0029,16'h0005,-16'h001d,16'h0010,16'h001d,16'h0024,16'h006e,-16'h00e0,16'h0043,16'h001b,-16'h002e,-16'h0001,16'h001c,16'h0002,-16'h0139,16'h000f,-16'h0019,16'h008f,16'h001e,-16'h0044,16'h004c,-16'h0097,16'h002d,16'h004b,-16'h0049,16'h0051,-16'h001a,16'h0052,16'h003b,16'h0057,-16'h0060,16'h000e,-16'h0049,16'h003b,16'h000d,-16'h005c,16'h0060,-16'h002b,16'h0024,16'h004e,16'h0083,16'h003b,16'h0057,-16'h006c,16'h0000,-16'h0025,16'h0068,-16'h0002,16'h0038,16'h006d,16'h006a,-16'h0022,16'h0031,16'h0040,16'h0010,16'h0053,-16'h0061,16'h0039,16'h006d,-16'h0023,16'h0013,-16'h000e,16'h000d,16'h008f,-16'h003d,16'h001b,16'h0001,16'h002f,16'h003d,16'h0051,16'h004b,-16'h005d,16'h0023,-16'h0021,-16'h0049,-16'h0049,16'h0017,-16'h0015,-16'h00f8,16'h000e,16'h001d,16'h0046,-16'h0020,-16'h0044,16'h003b,-16'h0077,16'h000d,16'h004f,-16'h003e,16'h005f,-16'h0007,16'h006a,16'h0036,16'h003f,-16'h0063,16'h0032,-16'h0030,-16'h0040,16'h0017,-16'h0085,16'h004c,16'h0023,-16'h0028,16'h0045,16'h007f,16'h0004,16'h0011,-16'h0062,16'h001e,-16'h005e,16'h0040,-16'h001f,16'h002a,16'h002c,16'h009a,16'h001c,16'h0033,16'h0071,-16'h001a,16'h003a,-16'h0077,16'h0035,16'h0051,-16'h000d,16'h0004,16'h000b,16'h0017,16'h0085,-16'h003a,-16'h0006,16'h0009,16'h0036,16'h003e,16'h0051,16'h003d,16'h005a,16'h0024,-16'h002c,-16'h0051,-16'h0026,16'h0019,-16'h0046,-16'h00d4,16'h0026,16'h0026,16'h0005,-16'h000c,-16'h0022,-16'h0018,-16'h00ad,16'h0003,16'h0051,16'h0039,16'h0019,16'h0019,16'h0098,16'h0064,16'h0023,16'h0016,16'h0029,-16'h0032,-16'h009a,16'h0012,-16'h0074,16'h003a,16'h0031,-16'h0068,16'h0046,16'h004c,-16'h0031,16'h0035,-16'h0072,16'h0043,-16'h0025,16'h0042,-16'h000a,16'h0034,16'h001e,16'h0092,16'h0061,16'h0029,16'h0078,16'h0006,16'h0034,-16'h0081,-16'h0008,16'h004c,-16'h002c,-16'h000e,16'h0027,-16'h0008,16'h0062,-16'h0017,-16'h0004,16'h000e,16'h002a,16'h0044,16'h0020,16'h004c,16'h00b6,16'h003f,-16'h0055,-16'h002e,-16'h001c,16'h0011,-16'h0044,-16'h00c3,16'h0017,16'h0041,-16'h000d,-16'h000c,-16'h0023,-16'h0074,-16'h008d,-16'h0016,16'h0057,16'h0036,-16'h002b,16'h0025,16'h005b,16'h0063,16'h0031,16'h0047,16'h000c,-16'h0016,-16'h009f,16'h0017,-16'h0080,16'h001e,16'h002f,-16'h00a4,16'h0045,16'h0039,-16'h0037,16'h001f,-16'h003f,16'h003a,-16'h000f,16'h0045,-16'h001e,16'h002d,-16'h0030,16'h008f,16'h006a,16'h002a,16'h004e,16'h0016,16'h0026,-16'h005d,16'h0039,16'h002a,-16'h0010,-16'h0005,16'h002d,-16'h0017,16'h0069,-16'h0004,-16'h0010,16'h003e,-16'h0003,16'h0022,16'h0051,16'h0027,16'h0092,16'h0032,-16'h0036,-16'h002e,-16'h0021,-16'h000d,-16'h0057,-16'h00a2,-16'h0016,16'h0006,16'h002b,-16'h0039,-16'h000f,-16'h00bd,-16'h0080,16'h0054,16'h0053,16'h004a,-16'h0046,16'h001d,16'h0000,16'h004b,16'h004e,16'h0057,-16'h001c,-16'h0025,16'h0005,16'h001a,-16'h0060,16'h0007,16'h0019,-16'h0054,16'h003f,16'h0043,16'h000b,16'h0036,-16'h0029,16'h001f,-16'h002a,16'h0041,-16'h0021,16'h000c,-16'h003e,16'h0063,16'h0049,16'h001f,16'h0055,16'h003c,16'h002d,-16'h0040,16'h003d,16'h0000,16'h0013,-16'h001c,16'h0044,16'h0012,16'h0060,16'h0001,-16'h0023,16'h0028,16'h0000,16'h000f,16'h0040,16'h000d,16'h009f,16'h000b,-16'h000e,-16'h0013,-16'h001a,-16'h0047,-16'h0060,-16'h0084,16'h0009,-16'h0004,16'h0038,-16'h0016,16'h0026,-16'h00bb,-16'h0057,16'h0042,16'h0064,16'h0046,-16'h004c,-16'h000e,-16'h0022,16'h0057,-16'h000c,16'h0072,-16'h004c,-16'h0023,16'h0020,16'h002b,-16'h0078,-16'h0002,-16'h000e,-16'h0052,16'h0025,16'h0039,-16'h000d,16'h001a,16'h0004,16'h001a,16'h0000,16'h0027,-16'h0022,16'h0000,-16'h005d,16'h0074,16'h0022,16'h000a,16'h0033,16'h0021,16'h0048,-16'h0016,16'h0039,-16'h0015,16'h001e,-16'h0016,16'h0061,16'h001a,16'h002e,16'h0013,-16'h001e,16'h0000,16'h0007,16'h003b,16'h0012,16'h0031,16'h008f,16'h001f,16'h000f,16'h000a,-16'h000e,-16'h0039,-16'h0061,-16'h0076,16'h0025,-16'h0007,16'h0014,-16'h0027,16'h000d,-16'h0057,-16'h0039,16'h0028,16'h0079,-16'h000a,-16'h0066,-16'h0007,-16'h0074,16'h005e,-16'h006c,16'h0071,-16'h0015,-16'h0012,-16'h0010,16'h0006,-16'h0074,16'h001b,-16'h0006,-16'h0038,16'h0019,16'h0079,-16'h0026,16'h0025,16'h0011,16'h0034,-16'h0018,16'h000a,-16'h0006,16'h0017,-16'h004e,16'h0059,-16'h003c,16'h0009,16'h000d,16'h0013,16'h0056,-16'h001f,16'h0034,-16'h0012,16'h0025,-16'h001e,16'h0041,16'h0017,16'h001f,16'h0015,-16'h003f,16'h0006,16'h000e,16'h0018,-16'h0014,16'h0013,16'h0055,16'h003d,16'h001c,16'h0006,-16'h000b,-16'h0010,-16'h007c,-16'h005d,16'h0019,-16'h0012,16'h000c,-16'h003f,-16'h0019,-16'h0021,-16'h0019,16'h005e,16'h008a,16'h0002,-16'h003f,-16'h000c,-16'h00ba,16'h004a,-16'h0091,16'h003c,16'h0000,16'h000a,16'h0012,16'h0006,-16'h005e,-16'h0007,16'h0028,-16'h0012,-16'h0014,16'h0045,-16'h0022,16'h0003,-16'h000d,16'h0033,16'h0000,16'h0025,16'h001b,-16'h0013,-16'h0029,16'h000a,-16'h008d,16'h001f,16'h001f,16'h0021,16'h0033,-16'h002b,16'h0040,-16'h0021,16'h0038,-16'h0003,16'h001c,16'h000c,16'h0021,16'h003c,-16'h0013,16'h002a,-16'h0012,16'h0013,-16'h0026,-16'h0021,16'h0036,16'h003f,16'h0027,16'h0018,16'h000f,-16'h0008,-16'h0078,-16'h0065,16'h0011,-16'h001c,-16'h004b,-16'h0007,-16'h000a,16'h000c,-16'h004a,16'h004f,16'h0094,-16'h000a,16'h0053,-16'h002a,-16'h0099,16'h0028,-16'h0085,16'h0016,-16'h0008,-16'h001e,16'h0002,16'h001d,-16'h001d,-16'h0012,16'h0011,16'h0034,-16'h0014,16'h001f,-16'h0013,16'h0001,16'h0003,16'h002e,16'h0003,16'h0034,16'h000a,-16'h0003,-16'h0033,-16'h0017,-16'h0050,16'h001f,16'h0023,16'h0016,16'h003e,-16'h0021,16'h0051,-16'h004f,16'h0054,-16'h0014,16'h0010,16'h0023,16'h003d,16'h002d,16'h001c,16'h0039,-16'h001d,16'h002b,16'h0003,-16'h001a,16'h0006,16'h0056,16'h0015,-16'h003a,-16'h0007,16'h0029,-16'h0060,-16'h005e,-16'h000d,-16'h0027,-16'h0031,16'h001a,-16'h0026,16'h001f,-16'h0036,16'h004b,16'h009d,-16'h0028,16'h004c,-16'h0002,-16'h008e,16'h0048,-16'h0013,16'h0024,16'h002a,16'h0011,16'h0029,16'h000b,-16'h0002,-16'h0008,16'h0006,16'h0040,-16'h0002,-16'h001e,-16'h0027,-16'h0001,16'h001c,16'h0037,-16'h0017,16'h0048,16'h0003,-16'h002a,-16'h0021,-16'h0034,16'h0002,16'h0015,16'h000a,16'h0000,16'h0056,-16'h0015,16'h0035,-16'h0048,16'h0022,-16'h0020,16'h001f,16'h0006,16'h0015,16'h0020,16'h0020,16'h002e,-16'h000c,16'h0034,16'h0017,16'h000b,-16'h0018,16'h0057,16'h0012,-16'h000f,16'h0004,16'h004a,-16'h006e,-16'h0040,-16'h0010,-16'h002b,16'h0008,16'h001c,-16'h0047,16'h004f,-16'h0023,16'h0007,16'h0072,-16'h0003,16'h0047,16'h0001,-16'h0078,16'h0052,16'h0050,-16'h0009,-16'h0019,-16'h001a,-16'h000a,16'h001a,16'h0011,16'h0004,16'h001b,16'h0065,16'h000f,-16'h000f,-16'h0005,16'h0003,16'h001e,16'h001e,16'h0001,16'h0043,16'h0014,-16'h002d,16'h0013,-16'h003f,-16'h000c,16'h0042,16'h000c,-16'h001c,16'h0064,-16'h0005,16'h003a,-16'h0061,16'h001f,-16'h0012,16'h000a,16'h0012,16'h003f,16'h001a,16'h0029,16'h0003,16'h000a,16'h0040,-16'h0003,16'h001c,-16'h0053,16'h0044,-16'h0020,-16'h000b,16'h0021,16'h0002,-16'h0065,-16'h0043,-16'h001c,-16'h0039,-16'h0004,16'h0011,-16'h001c,16'h0055,16'h000a,-16'h008c,16'h0067,16'h0025,16'h007a,16'h000e,-16'h002b,16'h0059,16'h0080,-16'h0019,-16'h004c,-16'h003d,-16'h0028,16'h0025,16'h003b,16'h0021,16'h003e,16'h0082,16'h0002,16'h0000,-16'h0018,16'h001a,16'h001d,16'h001d,-16'h001a,16'h003e,16'h0004,16'h0017,16'h0012,-16'h0035,-16'h000f,16'h0038,16'h0019,-16'h003d,16'h0074,16'h0036,16'h0052,-16'h001f,16'h0020,-16'h0048,16'h0006,16'h0002,16'h0024,16'h0002,16'h0052,16'h0008,16'h0035,16'h006a,16'h0002,16'h000d,-16'h002a,16'h003b,-16'h002b,16'h0000,16'h001a,-16'h001f,-16'h004f,-16'h0044,-16'h0049,-16'h003a,-16'h0005,16'h0026,-16'h0024,16'h0048,-16'h0022,-16'h0217,16'h0049,16'h0000,16'h0071,16'h0024,16'h0026,16'h0064,16'h005e,-16'h0040,-16'h004f,-16'h0023,-16'h0020,16'h0029,16'h0021,16'h002d,16'h0048,16'h0061,16'h0039,16'h0019,-16'h0017,16'h0057,16'h0010,16'h001c,-16'h0007,16'h0018,-16'h0010,-16'h0016,16'h0018,-16'h000b,-16'h0010,16'h003b,16'h0014,-16'h0064,16'h0078,16'h0022,16'h0053,-16'h000f,-16'h0011,-16'h003e,-16'h0004,16'h0001,16'h0015,-16'h000e,16'h001a,-16'h000f,16'h0050,16'h000d,16'h0002,16'h0051,16'h000d,16'h0013,-16'h000d,-16'h0055,16'h0001,-16'h0025,-16'h006e,-16'h0046,-16'h004a,-16'h00e3,16'h000a,16'h0057,-16'h0021,16'h004d,-16'h004f,-16'h028b,16'h0035,16'h0015,16'h0051,-16'h001b,16'h0055,16'h0033,-16'h0001,16'h000a,-16'h000b,-16'h000d,16'h0025,16'h0000,16'h000c,-16'h0002,16'h0039,16'h0037,16'h003c,16'h0026,-16'h000b,16'h003b,16'h001c,16'h0006,16'h001d,16'h0018,-16'h0010,-16'h000e,16'h002b,-16'h0012,16'h0024,16'h0048,-16'h0011,-16'h0046,-16'h001f,16'h003b,16'h004a,-16'h000d,-16'h001a,-16'h000d,-16'h0029,-16'h000f,16'h002d,-16'h006f,-16'h0029,-16'h0009,16'h003e,-16'h0033,16'h0026,16'h007c,16'h003b,16'h0024,16'h000b,-16'h009e,-16'h0017,-16'h004b,-16'h008b,-16'h0049,-16'h0020,-16'h012e,16'h0018,16'h0059,-16'h0012,-16'h000e,-16'h003b,-16'h0159,16'h0028,16'h000d,16'h001f,-16'h0083,16'h0057,16'h0051,-16'h0083,16'h002f,-16'h000b,-16'h000a,16'h005b,16'h0016,16'h0008,16'h0004,16'h001b,16'h0044,16'h0058,16'h0027,16'h000d,16'h004b,-16'h000d,16'h0013,16'h002b,16'h0013,-16'h0010,-16'h000f,16'h0018,16'h002b,16'h0060,16'h0040,16'h0017,-16'h002d,-16'h00ce,16'h0063,16'h003a,-16'h0075,16'h0008,-16'h000b,-16'h0035,-16'h0019,16'h0049,-16'h0064,-16'h004b,-16'h0023,16'h004a,-16'h00c1,16'h0053,16'h006c,16'h0054,16'h0035,16'h000f,-16'h004a,16'h0010,-16'h0016,-16'h007e,-16'h0044,-16'h001c,-16'h010e,16'h0018,16'h001d,-16'h0082,-16'h0048,-16'h0034,-16'h00d6,16'h002f,-16'h0038,-16'h00dd,-16'h0080,16'h007a,16'h002e,-16'h0107,16'h0049,16'h0018,-16'h0022,16'h0063,16'h000e,16'h0029,-16'h0013,-16'h0007,16'h004a,16'h005d,16'h0039,16'h0038,16'h0042,-16'h002a,-16'h0011,16'h0057,-16'h001c,-16'h0016,16'h0003,16'h001f,16'h002c,16'h0040,16'h0045,16'h000c,-16'h003d,-16'h00e3,16'h0066,16'h0033,-16'h005c,16'h0010,16'h0000,-16'h0036,-16'h0030,16'h0015,-16'h004e,-16'h003e,-16'h003b,16'h0026,-16'h00d6,16'h0071,16'h0054,16'h0074,16'h0031,16'h0027,-16'h003a,16'h0012,16'h0024,-16'h0071,-16'h0042,-16'h0012,-16'h00b2,-16'h0015,-16'h0054,-16'h00a4,-16'h0050,-16'h003e,-16'h0080,16'h0029,-16'h0028,-16'h01ce,-16'h0044,16'h002e,16'h003b,-16'h010d,16'h0042,16'h0052,-16'h002c,16'h0028,-16'h001c,16'h0052,-16'h0022,-16'h0001,16'h0070,16'h008b,16'h0058,16'h000e,16'h0048,-16'h0012,16'h0008,16'h0054,-16'h002b,16'h001d,-16'h001c,16'h000c,-16'h001b,16'h006b,16'h0026,16'h0024,-16'h002a,-16'h00a2,-16'h0017,16'h0060,-16'h005e,16'h0018,16'h0007,-16'h001a,-16'h002b,-16'h000a,-16'h0071,-16'h003c,-16'h0014,-16'h000c,-16'h00e9,16'h0034,16'h0033,16'h0071,16'h005c,16'h0015,16'h0009,16'h0008,-16'h0004,-16'h0074,-16'h0029,-16'h000b,-16'h006b,-16'h0042,-16'h0073,-16'h00d4,-16'h001e,-16'h001d,-16'h0038,16'h002a,-16'h000c,-16'h01a3,-16'h0015,-16'h0031,16'h0051,-16'h00c5,16'h003b,16'h0054,-16'h000e,16'h000b,-16'h001b,16'h0046,-16'h0031,-16'h0001,16'h0060,16'h0093,16'h0052,-16'h0019,16'h0023,-16'h0002,16'h0005,16'h0036,-16'h0007,-16'h0009,-16'h001d,-16'h0001,-16'h0015,16'h0058,16'h002e,-16'h0007,-16'h0031,-16'h002b,-16'h006a,16'h0047,-16'h0008,16'h005e,16'h0017,-16'h0031,-16'h002d,16'h001a,-16'h0052,-16'h0026,-16'h0017,-16'h0057,-16'h00c2,-16'h000e,-16'h0011,16'h0066,16'h0056,16'h0057,16'h0029,-16'h002c,-16'h002e,-16'h00b6,-16'h0018,16'h000e,-16'h0029,-16'h0087,-16'h0063,-16'h00b6,-16'h0029,-16'h000d,16'h0025,16'h0022,-16'h0009,-16'h013e,-16'h0024,-16'h0061,16'h007c,-16'h0072,16'h0030,16'h004c,16'h000b,-16'h0024,16'h0004,16'h0039,16'h0036,16'h000e,16'h002c,16'h008d,-16'h0010,-16'h0029,-16'h001b,-16'h002f,-16'h0028,16'h0011,16'h0013,-16'h0030,16'h000e,-16'h001b,-16'h004a,16'h000e,16'h0069,-16'h0034,-16'h002e,-16'h0007,-16'h00d6,16'h0078,-16'h006f,16'h0042,-16'h001c,16'h004f,16'h002a,16'h0000,16'h001f,16'h0029,16'h0052,16'h0024,16'h003c,-16'h0055,16'h0057,16'h005f,16'h0067,16'h004e,16'h0008,16'h0020,-16'h0056,16'h0021,-16'h0008,16'h0034,16'h000b,-16'h0016,16'h0066,16'h0020,16'h0016,-16'h00be,-16'h0066,16'h0013,-16'h005c,16'h004e,16'h00a0,16'h0030,16'h004a,16'h0013,-16'h000f,-16'h0017,16'h0017,-16'h0003,-16'h0009,16'h00ab,-16'h0002,16'h0027,16'h0043,16'h0038,16'h004a,-16'h0024,16'h001e,16'h000d,16'h0043,-16'h0036,-16'h0009,-16'h0001,-16'h0033,-16'h0034,-16'h00ac,16'h0030,-16'h0016,16'h0001,16'h001d,-16'h002b,-16'h0090,-16'h003a,-16'h0012,16'h0039,-16'h001a,16'h004a,16'h003a,16'h0031,-16'h0010,16'h0013,16'h0040,-16'h0008,16'h0031,-16'h0084,16'h0038,16'h001c,16'h0076,16'h0042,16'h0004,16'h0014,-16'h0029,16'h003c,-16'h0011,-16'h0012,16'h0008,-16'h003d,16'h0005,16'h0029,-16'h001e,-16'h0102,-16'h0041,-16'h000b,-16'h0070,16'h004e,16'h0076,16'h001d,16'h0065,16'h0026,-16'h0031,-16'h0027,-16'h0001,-16'h002b,-16'h0016,16'h00b7,16'h0046,16'h001a,16'h002b,16'h0053,16'h0052,-16'h0021,16'h000a,16'h0001,16'h0057,-16'h0041,-16'h002f,16'h0018,-16'h0031,16'h0023,-16'h00a4,16'h0050,-16'h0006,16'h0011,16'h0018,-16'h000b,-16'h0133,-16'h0030,16'h000e,16'h0032,-16'h0001,16'h0079,16'h002c,16'h0053,16'h000c,-16'h0004,16'h0020,16'h0001,16'h001d,-16'h0078,-16'h000a,-16'h0029,16'h0066,16'h000b,-16'h000d,16'h0000,-16'h000d,16'h0045,16'h001b,-16'h0021,16'h0018,-16'h0078,-16'h001c,16'h0058,-16'h007a,-16'h012d,-16'h0043,16'h000a,-16'h0073,16'h0001,16'h0050,16'h001f,16'h0031,16'h0023,16'h000e,-16'h001d,-16'h000b,-16'h0003,-16'h0006,16'h00a3,16'h001f,16'h001b,-16'h001c,16'h003f,16'h0062,-16'h002b,16'h001b,-16'h0030,16'h004f,16'h000a,-16'h0011,16'h0003,-16'h0025,16'h003d,-16'h0098,16'h0056,-16'h0014,16'h0003,16'h001f,16'h0004,-16'h016d,-16'h0021,16'h0029,16'h0017,16'h000a,16'h0072,16'h0024,16'h007b,16'h000f,-16'h0025,16'h0011,16'h0023,16'h0024,-16'h006a,-16'h0002,-16'h00ba,16'h004e,-16'h0066,16'h0001,-16'h0011,16'h002a,16'h0031,-16'h000d,-16'h003e,16'h0032,-16'h0082,-16'h004b,16'h0051,-16'h007f,-16'h014d,-16'h0026,16'h000b,-16'h0080,-16'h0011,16'h0074,-16'h000b,16'h002a,16'h001f,16'h004f,16'h0006,16'h0020,16'h0007,16'h001a,16'h0076,16'h0024,-16'h0008,-16'h0011,16'h003f,16'h0088,-16'h002e,-16'h001f,-16'h0062,16'h004b,16'h0027,16'h002f,16'h001b,-16'h0023,16'h0029,-16'h0074,16'h0070,-16'h0045,16'h0012,-16'h0001,16'h0055,-16'h0163,-16'h000b,16'h0023,16'h002b,16'h000b,16'h0072,16'h0029,16'h00c1,16'h0004,-16'h0055,16'h0011,16'h0036,16'h0020,-16'h0050,16'h002e,-16'h00fe,16'h0052,-16'h0073,16'h002c,-16'h0018,16'h0026,16'h0035,-16'h0026,-16'h0019,16'h003d,-16'h007d,-16'h0042,16'h00a9,-16'h0096,-16'h0112,-16'h0009,16'h0013,-16'h0019,-16'h002c,16'h003f,-16'h002c,-16'h0002,-16'h001b,16'h0085,16'h0026,-16'h0003,16'h0001,16'h0033,16'h0022,16'h000a,-16'h0018,-16'h0002,16'h003e,16'h0071,-16'h004c,-16'h0008,-16'h005b,16'h0018,16'h0008,16'h0084,16'h0004,-16'h002f,16'h0022,-16'h003f,16'h003e,-16'h0031,-16'h001f,-16'h0015,16'h005c,-16'h0199,16'h0005,16'h001b,16'h0020,16'h0008,16'h0044,16'h0004,16'h00a0,16'h000c,-16'h0045,-16'h0002,16'h0070,16'h0009,-16'h0038,16'h0040,-16'h00f4,16'h0065,-16'h0074,16'h0021,-16'h0004,-16'h0010,16'h003d,-16'h000d,-16'h0012,16'h0049,-16'h0048,-16'h0002,16'h00ab,-16'h0055,-16'h00ab,-16'h0003,16'h001e,16'h001b,-16'h0006,16'h0036,-16'h0087,-16'h001c,-16'h0043,16'h0084,16'h0035,-16'h0004,-16'h000a,16'h0033,16'h0021,-16'h0021,16'h0000,16'h0000,16'h0030,16'h0049,-16'h003f,-16'h001c,-16'h0048,16'h001c,16'h000a,16'h0091,16'h002a,-16'h0043,16'h003c,16'h000c,16'h0007,16'h0004,-16'h003c,-16'h0032,16'h0081,-16'h01b1,16'h0012,16'h0027,16'h0006,-16'h0001,16'h0036,16'h0002,16'h00ab,16'h001b,-16'h0047,16'h000b,16'h003a,16'h0027,-16'h0054,16'h004c,-16'h00ea,16'h006b,-16'h003a,16'h0052,16'h0007,-16'h0013,16'h0021,16'h001a,-16'h0016,16'h0022,-16'h001b,-16'h0005,16'h00af,16'h0047,-16'h00a0,16'h0013,16'h0025,16'h0040,16'h0029,16'h0047,-16'h009e,16'h0014,-16'h004b,16'h0090,16'h0021,-16'h0002,16'h0021,16'h0014,16'h0014,-16'h0031,-16'h0020,16'h001c,16'h0052,16'h005e,-16'h0041,16'h001c,-16'h0040,16'h0018,-16'h0013,16'h005e,-16'h000a,-16'h0036,16'h004b,16'h0019,-16'h0022,-16'h0002,-16'h0032,-16'h0015,16'h00a8,-16'h0176,16'h0013,16'h005b,16'h0003,16'h0019,16'h0031,16'h0008,16'h00c5,16'h001b,-16'h004e,16'h0010,16'h004a,16'h0023,-16'h0035,16'h0043,-16'h00c5,16'h007a,16'h0027,16'h003c,16'h0008,-16'h0012,16'h0045,16'h0018,-16'h002a,-16'h002a,16'h003d,16'h001a,16'h0089,16'h007a,-16'h00a6,16'h0032,16'h003a,16'h0000,16'h0042,16'h0031,-16'h0070,16'h0013,16'h0007,16'h0012,-16'h002e,-16'h000c,16'h005a,16'h0009,-16'h0012,-16'h005d,-16'h005f,16'h0042,16'h0041,16'h004f,-16'h000a,16'h004a,-16'h004d,16'h0023,-16'h0022,16'h006b,-16'h0008,-16'h0028,16'h0084,16'h0015,-16'h004a,16'h002f,-16'h0018,16'h0011,16'h008a,-16'h0166,16'h0027,16'h005d,-16'h0018,16'h0007,-16'h0009,16'h002c,16'h00b1,-16'h0008,-16'h003b,-16'h0013,16'h003a,16'h002c,16'h0000,16'h007f,-16'h00ab,16'h0071,16'h0026,16'h0021,-16'h000f,-16'h002a,16'h0045,-16'h000d,-16'h0018,-16'h003a,16'h006c,16'h0022,16'h0049,16'h005d,-16'h009b,16'h004f,16'h0048,-16'h0080,16'h0042,16'h0031,16'h0047,16'h002a,16'h003d,-16'h0029,-16'h0040,16'h000b,16'h0099,-16'h0002,-16'h0036,-16'h001c,-16'h0075,16'h0062,16'h005b,16'h0070,16'h001f,16'h0052,-16'h0032,16'h000b,-16'h0021,16'h0057,-16'h002f,16'h001e,16'h0073,16'h0064,-16'h0083,16'h0040,16'h0011,16'h0037,16'h008f,-16'h014a,16'h0020,16'h0046,-16'h0002,16'h000d,-16'h002c,16'h001b,16'h009f,-16'h002b,-16'h0023,16'h000c,16'h004e,16'h0032,16'h000e,16'h005b,-16'h0076,16'h004e,16'h0025,16'h0018,-16'h0032,-16'h001d,16'h004f,16'h001e,16'h0005,-16'h0018,16'h0069,16'h0012,16'h001b,16'h003f,-16'h0083,16'h0026,16'h006a,-16'h00ba,16'h0039,-16'h0015,16'h007a,16'h0035,16'h0044,-16'h005f,16'h0024,-16'h0003,16'h003b,-16'h000e,-16'h0033,16'h0074,-16'h002a,16'h0057,16'h0063,16'h009c,16'h0067,16'h0043,-16'h0040,16'h0023,-16'h0054,16'h0072,-16'h0027,16'h0002,16'h0032,16'h0071,-16'h0025,16'h0067,16'h003d,16'h002f,16'h00a1,-16'h00f3,16'h0038,16'h0054,16'h0008,16'h000e,-16'h001d,16'h001b,16'h0073,-16'h004f,-16'h0020,-16'h001e,16'h003c,16'h0051,16'h003d,16'h0030,16'h000f,16'h004c,-16'h0011,16'h0000,-16'h0022,-16'h0025,16'h0062,-16'h0003,16'h002d,16'h0022,16'h005e,16'h001d,16'h0002,-16'h0006,-16'h0088,16'h001e,16'h0049,-16'h004a,16'h003c,-16'h001e,16'h007b,16'h0046,16'h004e,-16'h0030,16'h0048,-16'h001c,-16'h004a,16'h0010,-16'h004d,16'h0058,16'h002f,16'h002e,16'h006c,16'h005e,16'h0050,16'h0017,-16'h004b,16'h0029,-16'h0051,16'h0084,-16'h0011,16'h0000,16'h0017,16'h0084,16'h003e,16'h004e,16'h0074,16'h001d,16'h00a2,-16'h00b2,16'h0019,16'h005b,-16'h000c,16'h000e,-16'h0010,-16'h0008,16'h008a,-16'h0043,-16'h0029,16'h0023,16'h002f,16'h0044,16'h002b,16'h0038,16'h0089,16'h0048,-16'h002d,-16'h0016,-16'h0015,-16'h0027,16'h0050,-16'h0022,16'h001f,16'h003d,16'h0018,-16'h0007,16'h0034,-16'h005a,-16'h0094,16'h0021,16'h0050,16'h0028,16'h0015,-16'h0009,16'h009b,16'h0030,16'h002c,16'h0020,16'h0000,-16'h0023,-16'h0080,-16'h0015,-16'h004b,16'h003f,16'h0049,-16'h0013,16'h0051,16'h003f,16'h0030,16'h001b,-16'h0039,16'h004c,-16'h002e,16'h004f,16'h0000,-16'h000b,16'h0005,16'h0078,16'h0064,16'h0058,16'h005e,16'h0029,16'h0085,-16'h008d,16'h0024,16'h0062,16'h0008,16'h0011,16'h0025,-16'h0029,16'h009b,-16'h0038,-16'h002b,16'h003b,16'h0029,16'h0009,16'h0041,16'h0031,16'h009b,16'h003b,-16'h004b,-16'h001a,-16'h001c,-16'h0035,16'h004c,-16'h0037,-16'h0007,16'h0059,16'h001c,-16'h0003,16'h001a,-16'h00a5,-16'h0099,-16'h001c,16'h004d,16'h0025,-16'h0018,16'h0011,16'h002b,16'h0021,16'h004d,16'h006d,-16'h002e,-16'h0011,-16'h0069,16'h000f,-16'h0030,16'h0039,16'h0068,-16'h0034,16'h0034,16'h0047,16'h0020,16'h002e,-16'h003c,16'h0019,-16'h0031,16'h0044,-16'h000a,-16'h0007,-16'h0024,16'h0073,16'h009a,16'h0058,16'h005e,16'h0035,16'h006d,-16'h0035,16'h002d,16'h0064,16'h0009,16'h0015,16'h0012,-16'h002b,16'h007a,16'h0000,-16'h0033,16'h0037,-16'h001d,-16'h0001,16'h0032,16'h0008,16'h0087,16'h0037,-16'h001e,-16'h001c,-16'h0033,-16'h0033,16'h0028,-16'h0049,-16'h0004,16'h0031,16'h0020,-16'h0020,16'h001d,-16'h00ac,-16'h0058,16'h0037,16'h0053,16'h000f,-16'h0033,16'h0033,-16'h0028,16'h0026,16'h0042,16'h0072,-16'h001c,-16'h001b,16'h0028,16'h002d,-16'h005c,-16'h0001,16'h001f,16'h001b,16'h0057,16'h0065,16'h0034,16'h002f,-16'h001c,16'h003d,-16'h0026,16'h003b,-16'h0013,-16'h0019,-16'h0033,16'h0078,16'h0070,16'h0047,16'h0053,16'h0036,16'h008e,-16'h0016,16'h003b,16'h0020,16'h000b,16'h0005,16'h002a,16'h000e,16'h005f,-16'h001f,-16'h002d,16'h0026,-16'h0037,16'h0006,16'h002e,16'h0027,16'h0087,16'h0033,-16'h000b,16'h0005,-16'h001b,-16'h0056,16'h003e,-16'h002a,16'h0010,16'h001b,16'h002e,-16'h001d,16'h0030,-16'h009d,-16'h002e,16'h004a,16'h002d,16'h0008,-16'h0064,16'h002f,-16'h007a,16'h003a,16'h0005,16'h0066,-16'h003c,-16'h0016,16'h0023,16'h0046,-16'h0068,16'h0027,16'h0002,16'h001f,16'h001d,16'h0053,16'h000d,16'h0021,16'h0013,16'h0020,-16'h0020,16'h0032,-16'h000e,-16'h002d,-16'h003a,16'h005a,16'h0017,16'h002a,16'h0054,16'h003d,16'h0086,-16'h0003,16'h0033,-16'h0007,16'h0022,-16'h0007,16'h0040,16'h001c,16'h0069,-16'h0012,-16'h0037,16'h001a,-16'h001f,16'h000a,16'h0002,16'h004a,16'h0071,16'h0060,16'h0015,16'h002a,-16'h002a,-16'h005b,16'h0038,-16'h004d,16'h000e,16'h0018,16'h0014,16'h0005,16'h0031,-16'h0077,-16'h0006,16'h003a,16'h0049,-16'h002c,-16'h007b,16'h0021,-16'h0079,16'h0035,-16'h0037,16'h0028,-16'h0025,16'h0005,16'h0033,16'h0034,-16'h005c,16'h0036,16'h000f,16'h0030,16'h0016,16'h0068,16'h000b,16'h0022,16'h0001,16'h001d,-16'h0010,16'h0028,16'h0003,-16'h0004,-16'h003c,16'h0055,-16'h0036,16'h0036,16'h003d,16'h002b,16'h007d,16'h000f,16'h003a,-16'h0011,16'h002d,16'h0019,16'h0045,16'h001f,16'h0050,16'h0021,-16'h0051,16'h0015,16'h0009,16'h0007,-16'h0040,16'h0048,16'h0056,16'h0066,16'h0012,16'h0021,16'h0003,-16'h002b,16'h002a,-16'h002a,16'h0020,16'h000c,-16'h0017,-16'h0022,-16'h0013,-16'h0025,-16'h0013,16'h006f,16'h005a,-16'h0025,-16'h003d,-16'h0012,-16'h0091,16'h0045,-16'h0068,16'h001e,-16'h0025,16'h0012,16'h002a,16'h0026,-16'h0050,16'h001a,-16'h0002,16'h0029,16'h0008,16'h0040,16'h000e,16'h0026,16'h000b,16'h0034,-16'h0019,16'h004e,16'h0018,-16'h0019,-16'h0023,16'h002c,-16'h009e,16'h0050,16'h0067,16'h001b,16'h0044,-16'h0004,16'h006a,-16'h0027,16'h0063,-16'h0003,16'h0029,16'h000f,16'h004c,16'h001a,-16'h0010,16'h0028,16'h000e,16'h000c,-16'h001a,16'h0000,16'h0046,16'h005f,16'h0009,-16'h0005,-16'h0002,-16'h0026,16'h004d,-16'h0029,16'h0004,16'h0017,-16'h003a,-16'h0014,-16'h003c,16'h0025,-16'h002b,16'h0062,16'h0071,-16'h0044,16'h005b,-16'h0054,-16'h0088,16'h002e,-16'h006c,16'h0000,16'h0008,16'h000f,-16'h0011,-16'h0007,-16'h0030,16'h0003,16'h0010,16'h002f,-16'h0008,16'h0041,-16'h0001,-16'h0013,16'h0026,16'h0031,-16'h001c,16'h0074,16'h000b,-16'h002b,-16'h0031,-16'h001b,-16'h004d,16'h0065,16'h0029,-16'h0002,16'h005c,-16'h001c,16'h0052,-16'h0047,16'h0041,16'h0003,16'h0029,16'h0008,16'h003d,16'h0022,16'h0002,16'h003b,-16'h0008,16'h0012,16'h0000,16'h0006,16'h0004,16'h0046,16'h001c,-16'h000d,-16'h0003,-16'h0008,16'h0010,-16'h0023,-16'h0012,-16'h0012,-16'h003e,16'h0019,-16'h0034,16'h004f,-16'h001f,16'h0062,16'h007c,-16'h0024,16'h0051,-16'h0034,-16'h0063,16'h002f,16'h000e,-16'h0015,16'h0026,16'h0022,-16'h001b,16'h0001,-16'h000a,16'h0000,16'h0045,16'h0039,16'h0031,-16'h0005,-16'h0004,-16'h0018,16'h0030,16'h0025,-16'h0009,16'h0055,16'h0008,-16'h0055,-16'h000c,-16'h0014,16'h003e,16'h0055,16'h002a,-16'h0013,16'h007f,-16'h0010,16'h003c,-16'h0059,16'h0037,-16'h0006,16'h0019,16'h001d,16'h0053,16'h0013,16'h003c,16'h002b,16'h0022,16'h0030,16'h000e,16'h0009,-16'h0014,16'h005e,-16'h0019,-16'h002a,16'h0008,-16'h0009,-16'h0005,-16'h0019,-16'h0026,16'h0000,16'h0002,16'h0018,-16'h0052,16'h0052,-16'h0039,16'h001f,16'h006f,16'h0010,16'h0063,-16'h0037,-16'h004e,16'h0040,16'h0051,-16'h000a,-16'h0021,-16'h0011,-16'h001a,16'h0004,16'h0017,16'h0003,16'h0034,16'h005f,16'h0005,16'h0015,16'h0003,-16'h000a,16'h001b,16'h001d,-16'h000d,16'h0044,16'h0005,-16'h0043,16'h0002,-16'h0020,16'h0036,16'h005b,16'h0022,-16'h0028,16'h0074,-16'h0021,16'h0041,-16'h0057,16'h001e,-16'h000e,-16'h001d,16'h002b,16'h0047,16'h002f,16'h004c,-16'h0015,16'h0023,16'h0027,-16'h002e,16'h0024,-16'h0053,16'h0041,-16'h000a,-16'h0003,16'h001b,-16'h0033,-16'h0015,-16'h001f,-16'h0034,16'h0029,-16'h000b,16'h0029,-16'h0036,16'h004f,-16'h0017,-16'h00ba,16'h0063,-16'h0029,16'h007d,-16'h002b,16'h0008,16'h0051,16'h007c,-16'h0004,-16'h004b,-16'h0026,-16'h002f,16'h0015,16'h0026,16'h001a,16'h0049,16'h0062,16'h0008,16'h000d,-16'h0011,-16'h0007,16'h000f,16'h0028,-16'h0013,16'h002f,-16'h0020,-16'h001f,16'h0023,-16'h0037,16'h0002,16'h004f,16'h0019,-16'h0026,16'h0092,16'h0012,16'h0039,-16'h003f,16'h0032,-16'h0043,-16'h002c,16'h003a,16'h003b,16'h001c,16'h0059,-16'h001d,16'h0043,16'h0012,-16'h0006,16'h003f,-16'h003a,16'h004a,-16'h000e,16'h0029,16'h001b,-16'h004a,-16'h001d,-16'h0033,-16'h0031,16'h0005,16'h0001,16'h006e,-16'h0012,16'h003d,-16'h002d,-16'h0228,16'h0059,-16'h0014,16'h003f,-16'h0012,16'h004b,16'h0034,16'h001e,-16'h0017,-16'h002e,-16'h0025,-16'h0007,16'h0024,16'h0017,16'h0043,16'h0059,16'h006a,16'h001f,16'h000e,-16'h0040,16'h001b,16'h000b,16'h001e,16'h0004,16'h0045,-16'h0015,-16'h0014,16'h000a,-16'h0011,16'h0013,16'h0057,16'h000b,-16'h001e,16'h007b,16'h004e,16'h002f,16'h0000,16'h0038,-16'h001d,-16'h002e,16'h000c,16'h0015,-16'h0005,16'h001a,-16'h002a,16'h0024,-16'h002d,16'h0013,16'h0059,16'h0006,16'h0039,-16'h0014,-16'h0031,16'h000d,-16'h0023,-16'h0032,-16'h0025,-16'h0036,-16'h0086,16'h002e,16'h0065,-16'h0032,16'h0024,-16'h005d,-16'h0294,16'h0057,-16'h001a,16'h0048,-16'h002d,16'h0060,16'h0027,-16'h000d,16'h0039,-16'h0014,-16'h001b,16'h0024,16'h0011,16'h0011,16'h0025,16'h004d,16'h0068,16'h0065,16'h0016,-16'h0033,16'h002a,16'h0022,16'h0008,16'h0000,16'h0038,-16'h0031,-16'h0028,16'h000d,-16'h001f,16'h003d,16'h0055,16'h0000,-16'h0011,-16'h002e,16'h001b,16'h0046,16'h0001,16'h0037,-16'h0027,-16'h0030,-16'h001a,16'h0031,-16'h0023,-16'h003f,-16'h0023,16'h004d,-16'h00e4,16'h0038,16'h0053,16'h0053,16'h0054,16'h000e,-16'h0035,16'h0005,-16'h0032,-16'h001b,-16'h002c,-16'h001f,-16'h00e1,16'h004c,16'h0041,-16'h005a,-16'h0015,-16'h0082,-16'h015f,16'h0048,-16'h000f,16'h0006,-16'h0053,16'h0062,16'h0026,-16'h0086,16'h004e,-16'h000c,-16'h000d,16'h0051,16'h0002,16'h0011,-16'h0006,16'h0002,16'h0056,16'h005e,16'h0016,-16'h000d,16'h0030,-16'h0012,16'h000c,16'h000b,16'h0017,-16'h0016,-16'h001d,16'h0041,-16'h001e,16'h005e,16'h006c,16'h0005,-16'h001c,-16'h0141,16'h003f,16'h002b,-16'h004d,-16'h0003,-16'h0011,-16'h003e,-16'h0038,16'h0038,-16'h003b,-16'h005c,-16'h0035,16'h0037,-16'h014c,16'h004b,16'h0058,16'h0052,16'h0050,16'h0001,-16'h0011,16'h0003,-16'h0013,-16'h004d,-16'h0030,16'h0000,-16'h00cc,16'h0022,-16'h0028,-16'h0089,-16'h0063,-16'h0039,-16'h00ce,16'h0054,-16'h0031,-16'h00d9,-16'h0065,16'h0057,16'h002f,-16'h00e4,16'h0052,16'h000f,-16'h0021,16'h003c,16'h0000,16'h0035,-16'h000e,-16'h0004,16'h0064,16'h008e,16'h003d,16'h0004,16'h0027,-16'h0007,16'h001f,16'h0042,-16'h0019,-16'h002f,16'h0008,16'h0027,-16'h0002,16'h003d,16'h005f,16'h0005,-16'h0021,-16'h014f,16'h005c,16'h001d,-16'h005a,16'h000c,16'h0009,-16'h000f,-16'h002a,16'h002d,-16'h0077,-16'h0035,-16'h002f,16'h0018,-16'h0192,16'h0058,16'h005e,16'h0065,16'h006c,16'h0006,-16'h0009,-16'h001f,-16'h0027,-16'h0047,-16'h0034,-16'h0011,-16'h00b0,-16'h0001,-16'h0098,-16'h00c0,-16'h0055,-16'h0046,-16'h0077,16'h0046,-16'h0019,-16'h01e7,-16'h002f,-16'h0003,16'h003d,-16'h00e9,16'h0052,16'h0049,-16'h0012,-16'h0009,-16'h0005,16'h0026,-16'h002c,-16'h001f,16'h008a,16'h00a2,16'h004c,-16'h004a,16'h003b,16'h0005,16'h002d,16'h004f,-16'h002b,-16'h0014,16'h0010,16'h000a,-16'h0017,16'h004f,16'h002f,16'h0011,-16'h0017,-16'h00c2,16'h0014,16'h002c,-16'h006e,16'h0010,16'h0021,16'h0008,-16'h0041,16'h0033,-16'h008f,-16'h0039,-16'h003a,-16'h000a,-16'h0144,16'h0028,16'h0051,16'h0065,16'h0035,16'h001e,16'h0009,-16'h0016,-16'h0016,-16'h004a,-16'h0024,-16'h0018,-16'h005e,-16'h0088,-16'h00a2,-16'h00c7,-16'h001a,-16'h0042,-16'h001f,16'h003c,-16'h0010,-16'h01b4,-16'h002d,-16'h002f,16'h0051,-16'h00aa,16'h0036,16'h0020,-16'h001d,-16'h0027,16'h0015,16'h003c,16'h0003,16'h0008,16'h006b,16'h00b3,16'h003a,-16'h003e,16'h0013,-16'h001e,16'h000b,16'h0042,-16'h0008,16'h000e,-16'h0021,16'h0011,-16'h000f,16'h0021,16'h0018,16'h0013,-16'h0013,-16'h0043,-16'h0048,16'h0032,-16'h0024,16'h004d,16'h000a,-16'h001e,-16'h0031,16'h0023,-16'h0096,-16'h001e,-16'h0036,-16'h004d,-16'h00f1,-16'h0004,16'h003d,16'h0050,16'h0047,16'h0035,16'h0029,-16'h005f,-16'h0015,-16'h0058,-16'h0021,16'h001d,-16'h0026,-16'h00ab,-16'h0097,-16'h00a4,-16'h0017,-16'h003b,16'h002e,16'h004c,16'h0000,-16'h011f,-16'h0023,-16'h0085,16'h005e,-16'h0063,16'h0011,16'h0023,16'h0028,-16'h0019,16'h0026,16'h0003,16'h0035,16'h001f,16'h0039,16'h00ad,-16'h002e,-16'h0079,-16'h0018,-16'h002c,-16'h0015,16'h002a,16'h0009,16'h0006,-16'h0003,16'h0003,-16'h002a,16'h0011,16'h0044,16'h0001,-16'h0014,-16'h0020,-16'h00c7,16'h0065,-16'h0038,16'h0068,16'h0003,16'h003c,16'h002d,-16'h0004,-16'h0013,16'h001d,16'h004e,16'h002f,16'h0040,-16'h0037,16'h00aa,-16'h0005,16'h0072,16'h004c,-16'h000f,16'h000e,-16'h0037,-16'h0015,-16'h0005,-16'h0010,-16'h0036,-16'h0011,16'h006f,16'h0021,-16'h0007,-16'h0092,-16'h003e,-16'h0010,-16'h0077,16'h002f,16'h00ac,16'h0023,16'h002f,16'h0020,-16'h002f,-16'h002b,16'h001b,16'h0000,-16'h0017,16'h0092,16'h0000,16'h0023,16'h0056,16'h0024,16'h0034,-16'h002d,16'h0007,16'h0001,16'h0045,-16'h002c,16'h0009,-16'h0009,-16'h0059,-16'h0009,-16'h0085,16'h002b,-16'h0008,-16'h001a,16'h0006,-16'h0037,-16'h005e,-16'h0043,-16'h0016,16'h0055,-16'h0008,16'h0037,16'h004e,16'h0009,-16'h0021,16'h0017,16'h002e,16'h0002,16'h001e,-16'h0049,16'h0047,-16'h0031,16'h007a,16'h0068,-16'h000d,16'h0015,-16'h0039,16'h0011,16'h0036,-16'h0024,16'h0012,-16'h0016,16'h0017,16'h003b,-16'h0041,-16'h00cd,-16'h0055,-16'h0012,-16'h009c,16'h003b,16'h0093,16'h001d,16'h004d,16'h002d,-16'h0039,-16'h0039,-16'h0006,16'h0019,-16'h0014,16'h008f,16'h0035,16'h0013,16'h002e,16'h0055,16'h004a,-16'h000d,16'h0020,16'h0004,16'h0035,-16'h0049,-16'h000f,-16'h0012,-16'h0014,16'h0031,-16'h007b,16'h0069,16'h0006,-16'h0006,16'h002b,-16'h0027,-16'h00bc,-16'h002e,16'h0006,16'h004f,16'h0014,16'h006c,16'h0060,16'h0031,-16'h000e,-16'h001d,16'h0024,16'h0003,16'h0011,-16'h003a,16'h0049,-16'h003c,16'h005c,16'h0026,-16'h0004,16'h000f,-16'h000c,16'h0033,16'h005c,-16'h0032,16'h0003,-16'h0062,-16'h0036,16'h005c,-16'h006e,-16'h0114,-16'h001a,-16'h001d,-16'h00a5,16'h0016,16'h005b,16'h001a,16'h0041,16'h0019,16'h0013,-16'h0035,16'h0001,16'h000c,16'h0017,16'h0066,16'h0036,16'h0000,16'h0008,16'h0050,16'h0033,-16'h001b,16'h000c,-16'h0008,16'h002b,16'h0009,-16'h0002,16'h0018,-16'h0034,16'h0022,-16'h0052,16'h0082,-16'h001f,16'h0011,16'h000f,16'h000f,-16'h0100,-16'h003c,16'h0025,16'h0020,16'h000a,16'h007a,16'h0030,16'h0053,-16'h001a,-16'h0013,16'h000e,16'h0016,16'h000f,-16'h0029,16'h000c,-16'h00ac,16'h003c,-16'h004a,-16'h0014,-16'h0020,16'h001c,16'h0030,16'h005e,-16'h0033,16'h001b,-16'h0059,-16'h0017,16'h0061,-16'h0077,-16'h0108,-16'h0027,16'h0002,-16'h00bb,-16'h0002,16'h004e,-16'h000e,16'h0019,-16'h0018,16'h0050,-16'h0014,-16'h000e,-16'h000b,16'h005b,16'h0050,16'h002a,-16'h0003,16'h0017,16'h004d,16'h0047,-16'h0023,-16'h0020,-16'h002d,16'h002a,-16'h0015,16'h0034,16'h0016,-16'h003f,16'h004d,16'h000e,16'h0062,-16'h004f,-16'h0013,-16'h0003,16'h0049,-16'h00fd,-16'h005a,16'h0014,16'h0041,16'h0006,16'h0067,16'h000e,16'h0064,-16'h001d,-16'h0042,16'h001a,16'h004b,16'h0007,-16'h0046,16'h0023,-16'h0110,16'h0045,-16'h006b,16'h0021,-16'h0013,16'h0005,16'h0044,16'h0076,-16'h000a,16'h0030,-16'h0076,16'h000f,16'h007b,-16'h004b,-16'h00f2,-16'h0008,-16'h000a,-16'h0056,16'h000a,16'h005f,16'h0014,16'h0000,-16'h0032,16'h008c,16'h0000,16'h0016,-16'h002e,16'h0050,16'h001e,16'h0015,-16'h001a,16'h0013,16'h0055,16'h0061,-16'h003a,-16'h0005,16'h000a,16'h001a,16'h0019,16'h0063,16'h0015,-16'h0045,16'h0038,16'h0046,16'h0055,-16'h000d,-16'h001b,-16'h0034,16'h005d,-16'h0129,-16'h003a,16'h000b,16'h0046,16'h0011,16'h004e,16'h001f,16'h0081,-16'h000a,-16'h003f,-16'h000c,16'h0070,16'h0010,-16'h0038,16'h003f,-16'h0154,16'h006f,-16'h0058,16'h001a,-16'h0016,16'h0003,16'h0031,16'h0082,-16'h0004,16'h0041,-16'h0057,-16'h0001,16'h00af,16'h000b,-16'h00a4,16'h0002,16'h001c,-16'h0005,16'h0003,16'h003d,-16'h0027,-16'h0015,-16'h006b,16'h0089,16'h0020,-16'h0003,-16'h0021,16'h0042,-16'h000e,-16'h0013,16'h000a,-16'h0015,16'h0081,16'h0042,-16'h0050,16'h0024,16'h001e,-16'h000e,16'h001c,16'h006a,16'h0013,-16'h0041,16'h003c,16'h0044,16'h002c,-16'h000b,-16'h0040,-16'h003c,16'h0062,-16'h0125,-16'h0021,16'h002d,16'h002c,16'h001a,16'h0043,16'h001c,16'h0090,-16'h0011,-16'h0021,16'h000d,16'h007d,16'h0012,-16'h0033,16'h0030,-16'h00d8,16'h005f,-16'h0025,16'h0013,-16'h0031,-16'h001c,16'h002f,16'h0088,16'h0000,16'h0057,16'h0003,16'h000e,16'h00d9,16'h0097,-16'h009d,16'h0014,16'h0020,-16'h000c,16'h001e,16'h0059,-16'h0028,16'h0011,-16'h0041,16'h0082,-16'h0038,-16'h0015,-16'h000a,16'h0026,-16'h0011,-16'h0032,-16'h0016,-16'h0008,16'h0069,16'h003e,-16'h0027,16'h003a,16'h001d,16'h0000,16'h0009,16'h006f,16'h0004,-16'h003e,16'h0030,16'h003e,-16'h001d,16'h0004,-16'h004e,-16'h0030,16'h0080,-16'h0116,-16'h0019,16'h001c,16'h004e,16'h000d,16'h0023,16'h0027,16'h005c,-16'h0004,-16'h001d,16'h0020,16'h0085,16'h0026,-16'h003d,16'h004a,-16'h00ae,16'h0077,16'h0027,16'h0024,16'h0000,16'h0001,16'h001f,16'h0099,-16'h000f,-16'h0019,16'h0022,16'h0020,16'h0099,16'h00aa,-16'h00a3,16'h0030,16'h0036,-16'h0081,16'h0018,16'h006a,16'h0011,16'h0025,16'h0018,16'h0017,-16'h0046,-16'h0013,16'h005c,16'h000c,-16'h002f,-16'h0036,-16'h006f,16'h0026,16'h006b,16'h0047,-16'h0017,16'h0059,16'h0016,16'h002b,-16'h0018,16'h008e,16'h0004,-16'h0037,16'h003c,16'h0069,-16'h0057,16'h0023,-16'h0032,16'h002f,16'h0068,-16'h010f,-16'h0018,-16'h0008,16'h0028,16'h0011,16'h000b,16'h000c,16'h0080,-16'h0010,-16'h002f,16'h0038,16'h0061,16'h0036,-16'h002a,16'h0071,-16'h006e,16'h0076,16'h0018,16'h0047,-16'h000c,-16'h0023,16'h0027,16'h0082,16'h0008,-16'h0014,16'h004f,16'h0058,16'h0086,16'h0056,-16'h0083,16'h0028,16'h0046,-16'h00e3,16'h0029,16'h001a,16'h0069,16'h003b,16'h001d,-16'h004e,-16'h001d,-16'h000b,16'h007e,16'h002c,-16'h0046,16'h0020,-16'h0099,16'h003a,16'h006c,16'h0065,16'h0009,16'h0038,16'h0021,16'h0037,-16'h0034,16'h009d,-16'h0025,-16'h002a,16'h0038,16'h0083,-16'h007f,16'h0043,-16'h0022,16'h004c,16'h0083,-16'h00d2,-16'h000e,-16'h000b,16'h0042,16'h000b,-16'h001c,16'h0014,16'h0061,-16'h001d,-16'h0003,16'h0020,16'h0073,16'h0039,-16'h0025,16'h0041,-16'h001d,16'h005b,16'h0006,16'h0073,-16'h0003,-16'h0033,16'h0038,16'h0072,16'h0023,16'h0013,16'h007d,16'h0032,16'h0042,16'h003b,-16'h007c,16'h0020,16'h0060,-16'h00d3,16'h0023,-16'h0027,16'h0085,16'h0046,16'h0023,-16'h004c,16'h0043,-16'h0014,16'h0003,16'h000f,-16'h002e,16'h006f,-16'h0062,16'h0029,16'h0089,16'h0063,16'h0028,16'h0026,16'h0018,16'h0018,-16'h0068,16'h009b,-16'h0013,-16'h0038,-16'h001d,16'h004c,-16'h0034,16'h002f,16'h0021,16'h003b,16'h0098,-16'h0081,-16'h0014,16'h0001,16'h0042,16'h001b,-16'h000a,16'h0027,16'h0071,-16'h0028,-16'h001a,16'h0030,16'h0063,16'h0028,-16'h0006,16'h0007,16'h0056,16'h005c,16'h0000,16'h004d,-16'h000a,-16'h0042,16'h0048,16'h0072,16'h0030,-16'h0008,16'h0068,16'h003b,16'h0048,-16'h0045,-16'h006f,16'h001b,16'h005a,-16'h0039,16'h0021,-16'h0054,16'h0099,16'h0031,16'h002a,-16'h0011,16'h0059,16'h0000,-16'h007b,-16'h000a,-16'h0035,16'h0041,16'h0029,16'h0018,16'h0079,16'h0044,16'h002c,16'h0002,16'h000c,16'h0020,-16'h008b,16'h0094,-16'h0001,-16'h0022,-16'h000a,16'h0046,16'h0025,16'h004f,16'h0053,16'h002f,16'h009b,-16'h006f,-16'h0009,16'h001f,16'h0023,16'h0000,16'h0007,16'h001e,16'h006e,16'h0004,-16'h0017,16'h0035,16'h0040,16'h001a,-16'h000a,16'h004c,16'h009c,16'h004f,-16'h0039,16'h0013,-16'h001a,-16'h004a,16'h004b,16'h0059,16'h002c,16'h0018,16'h003d,16'h0009,16'h0057,-16'h0086,-16'h0055,-16'h000f,16'h0037,16'h0021,16'h0021,-16'h0056,16'h0061,16'h0026,16'h003d,16'h001a,16'h0018,-16'h0014,-16'h008d,16'h0016,-16'h0004,16'h002c,16'h0040,16'h0020,16'h0059,16'h0048,16'h0040,16'h001e,-16'h0004,16'h000e,-16'h0040,16'h007e,16'h0027,-16'h004b,-16'h002e,16'h0020,16'h004e,16'h004f,16'h0036,16'h0032,16'h0084,-16'h0068,16'h0009,16'h001b,16'h0029,16'h000d,16'h0027,-16'h0011,16'h007f,16'h001c,-16'h003a,16'h0027,16'h0049,-16'h001c,16'h0014,16'h0014,16'h0085,16'h0028,-16'h002d,-16'h0005,-16'h0022,-16'h002d,16'h0052,16'h004d,-16'h0004,16'h002f,16'h002b,-16'h0035,16'h0028,-16'h00ad,-16'h0083,-16'h003b,16'h0054,16'h0015,-16'h001c,-16'h0010,16'h000d,16'h001c,16'h005a,16'h0079,-16'h0014,-16'h0014,-16'h0069,16'h000e,16'h000d,16'h000d,16'h0038,16'h0005,16'h0047,16'h0033,16'h003b,16'h0023,16'h0006,16'h002c,-16'h001f,16'h006b,16'h002a,-16'h0031,-16'h0044,16'h0035,16'h0088,16'h0041,16'h0046,16'h0047,16'h0081,-16'h001f,16'h002a,16'h0021,16'h0039,16'h0004,16'h001a,16'h0001,16'h0072,16'h0009,-16'h001b,16'h0037,16'h0017,-16'h0032,16'h000d,-16'h001b,16'h0066,16'h0039,-16'h0018,-16'h001f,-16'h001c,-16'h003a,16'h0055,16'h001c,16'h0013,16'h0022,16'h000f,-16'h003f,16'h0044,-16'h00a5,-16'h0061,16'h0040,16'h003d,16'h0002,-16'h0041,16'h0030,-16'h0046,16'h0020,16'h003d,16'h007b,-16'h0032,-16'h0004,16'h0046,16'h0005,-16'h0006,16'h0003,16'h0034,16'h0041,16'h0030,16'h004f,16'h004a,16'h0025,-16'h0005,16'h0023,-16'h0012,16'h003e,16'h0004,-16'h002b,-16'h000b,16'h001c,16'h008d,16'h0049,16'h0068,16'h003a,16'h0083,16'h0010,16'h002f,16'h0006,16'h0026,16'h0023,16'h0032,16'h0011,16'h0045,16'h0014,-16'h0019,16'h0012,-16'h0008,16'h0000,16'h001b,16'h0013,16'h0072,16'h003f,16'h0006,-16'h0008,-16'h0018,-16'h0051,16'h004f,16'h001f,16'h002c,16'h0026,16'h0020,16'h0003,16'h0070,-16'h008e,-16'h0011,16'h007d,16'h0043,-16'h0007,-16'h004d,16'h0054,-16'h00b6,16'h002d,16'h0017,16'h006e,-16'h001c,-16'h001f,16'h004c,16'h0020,-16'h001e,16'h004b,-16'h0001,16'h0061,16'h0023,16'h002a,16'h0022,16'h003c,16'h000b,16'h0014,-16'h000d,16'h004c,-16'h0013,-16'h0044,-16'h003c,16'h002d,-16'h001c,16'h0034,16'h007b,16'h0019,16'h008a,16'h003d,16'h003b,-16'h000d,16'h0026,16'h0019,16'h005b,16'h003a,16'h0046,16'h0008,-16'h0026,16'h0005,-16'h000b,16'h0007,-16'h000a,16'h003e,16'h006d,16'h0028,16'h000c,16'h000c,-16'h0011,-16'h0057,16'h0063,16'h001d,16'h0005,16'h002a,-16'h000c,16'h0006,16'h0076,-16'h0011,16'h001a,16'h0065,16'h0051,-16'h002f,-16'h0066,16'h0040,-16'h008d,16'h0029,16'h0024,16'h002c,16'h0010,16'h0002,16'h002d,16'h0046,-16'h002e,16'h002e,16'h002e,16'h0050,16'h003b,16'h0047,16'h002f,16'h0038,16'h001a,16'h0012,-16'h0025,16'h0066,-16'h0002,-16'h0018,-16'h0039,16'h0034,-16'h0063,16'h004b,16'h006d,16'h002e,16'h0096,16'h0054,16'h0047,16'h000b,16'h0028,16'h002c,16'h0059,16'h001e,16'h0025,16'h0018,-16'h0042,16'h000a,-16'h0003,-16'h000e,16'h0000,16'h0040,16'h0052,16'h003a,16'h0007,16'h0013,16'h0005,-16'h0047,16'h0083,16'h0014,-16'h0007,16'h0012,-16'h000e,16'h0012,16'h001c,16'h001f,16'h0000,16'h0084,16'h0048,-16'h004f,-16'h003e,16'h000b,-16'h008b,16'h0025,-16'h000f,16'h0017,16'h0012,16'h0018,16'h0030,16'h000d,-16'h0062,16'h000a,16'h0017,16'h004c,16'h001f,16'h003e,16'h000b,16'h000e,16'h000e,16'h002e,16'h0027,16'h0076,16'h0002,-16'h0008,-16'h0008,16'h0012,-16'h0091,16'h004b,16'h0075,16'h001c,16'h006e,16'h0030,16'h004b,-16'h0034,16'h0040,16'h0007,16'h0050,16'h002b,16'h0048,16'h000a,16'h0013,16'h0043,-16'h0001,16'h0003,16'h000d,16'h0004,16'h0039,16'h0030,16'h0010,16'h0030,-16'h0005,-16'h0040,16'h009e,16'h0023,-16'h0005,16'h0031,-16'h0030,16'h0010,-16'h0006,16'h003e,-16'h0022,16'h0086,16'h0055,-16'h003e,16'h003b,-16'h0033,-16'h009a,16'h0006,-16'h001e,-16'h0009,16'h0025,16'h0023,-16'h0016,-16'h0010,-16'h005f,16'h0004,16'h001d,16'h0048,16'h0020,16'h0032,16'h0009,-16'h0016,16'h0004,16'h0042,16'h0021,16'h007b,16'h0008,-16'h0019,16'h0004,16'h000e,-16'h004f,16'h0071,16'h0059,16'h0011,16'h0072,16'h0043,16'h004f,-16'h0061,16'h003f,16'h001f,16'h000c,16'h0019,16'h003b,16'h0002,16'h003c,16'h0029,16'h0021,-16'h000c,16'h0045,-16'h0003,16'h0015,16'h0029,-16'h0004,16'h000a,-16'h000f,-16'h0025,16'h0084,16'h002d,-16'h0018,16'h0029,-16'h002f,16'h001b,-16'h0040,16'h004d,16'h0004,16'h0059,16'h007b,-16'h0025,16'h0063,-16'h0038,-16'h003b,16'h0009,16'h002a,-16'h0025,16'h001b,16'h002b,-16'h0026,-16'h000e,-16'h003f,16'h0019,16'h006c,16'h0050,16'h002d,16'h003a,16'h0024,-16'h0001,16'h001d,16'h000b,16'h0014,16'h0065,-16'h0019,-16'h0048,-16'h000f,16'h000e,16'h001b,16'h0051,16'h0048,16'h000e,16'h0081,16'h0022,16'h0043,-16'h0052,16'h004c,16'h0010,16'h0022,-16'h0005,16'h003f,16'h0012,16'h0043,-16'h0009,16'h003d,-16'h002e,16'h000e,16'h0014,16'h0002,16'h0024,-16'h000c,16'h0011,16'h0032,-16'h0017,16'h005e,16'h002e,-16'h0004,16'h001f,-16'h0021,16'h002a,-16'h002a,16'h0053,-16'h0022,16'h0034,16'h006f,-16'h0021,16'h006d,-16'h002f,-16'h001e,16'h0004,16'h0032,-16'h0018,-16'h0015,16'h000d,-16'h000b,-16'h0001,-16'h001c,16'h0017,16'h0036,16'h0036,16'h0048,16'h003d,16'h002f,-16'h0009,16'h001c,16'h000a,16'h0001,16'h0073,-16'h0001,-16'h0034,-16'h0007,16'h0003,16'h0032,16'h003b,16'h0040,-16'h0004,16'h0097,-16'h0002,16'h0022,-16'h0062,16'h0023,16'h0009,-16'h0007,16'h0017,16'h0044,16'h0036,16'h0047,-16'h0021,16'h0029,-16'h0014,16'h0006,16'h0019,-16'h002b,16'h0031,-16'h002a,16'h001e,16'h0027,-16'h0035,16'h0050,16'h0015,-16'h0015,16'h0060,16'h0011,16'h0031,-16'h002d,16'h003c,-16'h0008,-16'h00b6,16'h0064,-16'h004c,16'h007f,-16'h0032,16'h0027,16'h0044,16'h0059,-16'h0015,-16'h0033,16'h0015,-16'h0020,-16'h0016,-16'h0004,16'h0024,16'h0035,16'h0038,16'h001c,16'h0048,16'h0000,16'h0012,-16'h0010,16'h0029,-16'h0002,16'h0040,-16'h0031,-16'h0018,16'h000e,-16'h0026,16'h0012,16'h0041,16'h0031,-16'h0027,16'h0099,16'h000d,16'h0006,-16'h001e,16'h0055,-16'h0023,-16'h001d,16'h0024,16'h0035,16'h0023,16'h0054,-16'h0027,16'h0022,-16'h005b,-16'h0009,16'h0041,-16'h0051,16'h004e,16'h0012,16'h001c,16'h0018,-16'h0029,16'h005b,16'h0005,-16'h0008,16'h003c,16'h0025,16'h0050,-16'h0040,16'h0037,-16'h0055,-16'h0248,16'h0034,-16'h0038,16'h0064,-16'h000d,16'h0031,16'h0017,16'h002a,16'h0027,-16'h0030,-16'h0009,-16'h0014,-16'h000f,16'h0039,16'h0039,16'h0034,16'h0050,16'h0026,16'h002c,-16'h0039,-16'h000c,16'h000d,16'h0041,16'h000e,16'h004e,-16'h0023,-16'h0032,16'h0008,-16'h0029,16'h002f,16'h0036,16'h000d,-16'h0015,16'h0056,16'h001c,16'h0011,16'h0009,16'h0047,-16'h0027,-16'h003d,16'h0002,16'h0023,16'h0027,-16'h0004,-16'h0034,16'h0018,-16'h00fd,16'h0021,16'h003c,16'h001a,16'h003f,-16'h0005,-16'h000b,16'h0001,-16'h002d,16'h0026,-16'h0005,16'h0001,-16'h003b,16'h003d,16'h0038,-16'h004c,16'h0027,-16'h0076,-16'h028f,16'h0059,-16'h0033,16'h005c,-16'h000b,16'h0047,16'h0009,16'h0000,16'h0042,-16'h0012,-16'h0005,-16'h0002,-16'h0014,16'h003c,16'h0023,16'h0056,16'h0070,16'h004c,16'h0012,-16'h0038,16'h0007,16'h0011,16'h0011,16'h000a,16'h005c,-16'h002d,-16'h0044,-16'h0005,-16'h0064,16'h003b,16'h0053,16'h0002,16'h0000,-16'h0090,16'h0018,16'h0031,16'h0002,16'h002b,-16'h002c,-16'h0022,-16'h001f,16'h0039,-16'h0001,-16'h001e,-16'h0043,16'h003a,-16'h017c,16'h0033,16'h004c,16'h0042,16'h0034,16'h000a,16'h0000,16'h0006,-16'h002c,16'h003b,-16'h0011,-16'h0006,-16'h00cb,16'h004f,-16'h0016,-16'h006c,-16'h0031,-16'h0055,-16'h0164,16'h0038,-16'h001b,16'h0026,-16'h003c,16'h0056,16'h0012,-16'h005c,16'h006a,-16'h000a,-16'h0021,16'h0046,-16'h0015,16'h0028,16'h0030,16'h0017,16'h003f,16'h004e,16'h0024,-16'h0013,16'h0032,16'h0000,16'h000d,-16'h0015,16'h0055,-16'h002c,16'h0001,16'h000a,-16'h0041,16'h0052,16'h004d,-16'h0006,16'h0016,-16'h01b5,16'h002f,16'h0016,-16'h0023,16'h0004,-16'h0017,-16'h0036,-16'h0030,16'h003e,16'h0009,-16'h0049,-16'h0044,16'h004c,-16'h01c4,16'h0053,16'h006c,16'h006a,16'h0036,16'h002c,16'h0012,16'h000e,-16'h0046,16'h002d,16'h000c,16'h0006,-16'h00b6,16'h0034,-16'h0082,-16'h0081,-16'h0071,-16'h002a,-16'h00e0,16'h004c,-16'h0027,-16'h00e0,-16'h004e,16'h0026,16'h0022,-16'h00a2,16'h0054,16'h0029,-16'h0021,16'h0030,-16'h0012,16'h002c,-16'h0005,-16'h0004,16'h0064,16'h0086,16'h002a,-16'h0033,16'h0042,16'h0015,16'h0020,16'h002e,-16'h0006,-16'h0002,16'h0017,-16'h001d,16'h0007,16'h0039,16'h004d,16'h0000,16'h0000,-16'h01bb,16'h0055,16'h001c,-16'h0043,16'h0008,-16'h0002,16'h0002,-16'h0048,16'h0028,-16'h0036,-16'h002c,-16'h0039,16'h002b,-16'h0159,16'h0059,16'h006a,16'h006f,16'h0028,16'h0004,-16'h000f,-16'h001b,-16'h001f,16'h0017,-16'h0009,-16'h000f,-16'h008d,-16'h0030,-16'h00af,-16'h0092,-16'h002f,-16'h0064,-16'h0069,16'h005d,-16'h001f,-16'h01d9,-16'h0031,-16'h001a,16'h001c,-16'h0082,16'h0043,16'h003c,16'h0016,16'h000e,-16'h0009,16'h0023,16'h000b,-16'h0010,16'h0092,16'h008b,16'h0021,-16'h003b,16'h002d,-16'h0002,16'h0022,16'h004b,16'h0000,-16'h001a,-16'h0008,16'h0017,16'h0008,16'h001c,16'h0039,16'h0026,-16'h0002,-16'h00f1,-16'h000f,16'h002c,-16'h006a,16'h004c,16'h0008,16'h0018,-16'h004b,16'h0047,-16'h008d,-16'h000d,-16'h0037,-16'h001b,-16'h011b,16'h004d,16'h005e,16'h005c,16'h002f,16'h0026,16'h0003,-16'h0044,-16'h0009,16'h0000,-16'h0002,-16'h0005,-16'h0040,-16'h007a,-16'h00c7,-16'h00ad,16'h0004,-16'h0046,-16'h000e,16'h004d,-16'h0007,-16'h01a0,16'h0000,-16'h0072,16'h0017,-16'h0059,16'h001b,16'h0032,16'h0009,16'h0014,16'h000f,16'h000d,16'h0005,-16'h0015,16'h009b,16'h008a,16'h001e,-16'h0069,16'h000f,-16'h0016,16'h0005,16'h0047,-16'h000c,16'h0019,16'h0014,16'h002b,16'h0003,16'h0010,16'h0027,16'h003a,16'h002a,-16'h006e,-16'h0046,16'h001c,-16'h0019,16'h003b,-16'h0008,16'h001a,-16'h0040,16'h0023,-16'h00b3,-16'h0005,-16'h004d,-16'h004d,-16'h00ed,16'h0000,16'h0033,16'h004d,16'h0024,16'h0038,16'h0031,-16'h0064,-16'h000e,16'h0008,-16'h000e,16'h0002,-16'h0007,-16'h008d,-16'h0087,-16'h0077,-16'h001e,-16'h0035,16'h002f,16'h0075,16'h0020,-16'h0111,16'h0004,-16'h0098,16'h0065,-16'h0032,16'h0004,16'h0010,16'h001f,16'h000a,16'h002d,16'h0017,16'h0026,16'h0028,16'h0074,16'h00bf,-16'h0031,-16'h0085,-16'h0029,-16'h0033,-16'h0017,16'h0055,16'h0014,16'h0017,-16'h0001,16'h0020,-16'h0027,16'h0012,16'h0038,16'h0002,16'h0012,-16'h004a,-16'h0085,16'h0035,-16'h000b,16'h005e,16'h0009,16'h0059,16'h004c,-16'h0009,16'h0003,16'h0035,16'h0046,16'h0031,16'h0048,-16'h002d,16'h00bb,-16'h0037,16'h0071,16'h0033,16'h0000,16'h001a,-16'h0021,-16'h0029,16'h0000,-16'h0006,-16'h0037,16'h000e,16'h0093,-16'h0002,16'h0000,-16'h00a0,-16'h006b,16'h0002,-16'h0042,16'h0029,16'h00d2,16'h0065,16'h0030,16'h003c,-16'h0042,-16'h0037,-16'h0003,-16'h0010,-16'h001a,16'h00ab,-16'h0020,16'h001a,16'h0063,16'h002c,16'h0003,-16'h0004,16'h000f,16'h0006,16'h0043,-16'h004b,16'h0013,-16'h0008,-16'h0030,16'h0037,-16'h0077,16'h0026,16'h000e,-16'h0046,-16'h0001,-16'h0025,-16'h002a,-16'h0040,16'h0032,16'h0047,16'h0003,16'h005a,16'h0066,16'h000d,-16'h003b,16'h002d,16'h0024,16'h001c,16'h0035,16'h0009,16'h0087,-16'h004a,16'h007c,16'h0034,16'h0014,16'h0013,-16'h002e,16'h0006,16'h001f,-16'h0029,-16'h0010,-16'h001f,16'h000b,16'h004b,-16'h0036,-16'h00d0,-16'h002c,-16'h002c,-16'h0064,16'h001e,16'h0071,16'h0041,16'h0043,16'h0043,-16'h0042,-16'h0030,-16'h0022,-16'h0001,16'h0006,16'h008f,16'h000f,16'h0009,16'h0053,16'h0054,16'h001d,16'h0002,16'h0026,-16'h0014,16'h002c,-16'h003b,-16'h0005,-16'h000a,-16'h0010,16'h0028,-16'h0056,16'h0047,-16'h0014,-16'h0006,16'h000d,-16'h002a,-16'h0077,-16'h004f,16'h0017,16'h004d,16'h0021,16'h0064,16'h0074,-16'h0015,-16'h003e,16'h0014,16'h002c,-16'h0002,16'h0016,16'h0024,16'h005b,-16'h0068,16'h006d,16'h0008,16'h0016,16'h000b,16'h0000,16'h0027,16'h0054,-16'h0022,-16'h0002,-16'h004d,-16'h0030,16'h0057,-16'h0053,-16'h0105,-16'h001c,-16'h0035,-16'h0094,16'h000c,16'h005b,16'h0017,16'h002e,16'h001c,-16'h0001,-16'h001f,-16'h0026,-16'h0016,16'h002d,16'h0061,16'h0030,-16'h000d,16'h002f,16'h005c,16'h003c,16'h0013,16'h0018,16'h000d,16'h0014,-16'h002e,16'h0005,-16'h0005,-16'h0027,16'h003f,-16'h0006,16'h0063,-16'h0012,16'h0001,-16'h001d,-16'h001a,-16'h007a,-16'h0068,-16'h0003,16'h002c,16'h000d,16'h0067,16'h004e,-16'h0011,-16'h001f,-16'h0003,16'h0005,-16'h001a,16'h0019,16'h0001,16'h000b,-16'h00ab,16'h0051,-16'h0015,16'h000b,-16'h0001,16'h0007,16'h002f,16'h005e,-16'h0043,16'h0000,-16'h0079,-16'h001a,16'h005a,-16'h0044,-16'h010e,-16'h001f,-16'h002e,-16'h005c,-16'h001c,16'h0042,-16'h001f,16'h001d,-16'h0025,16'h0041,-16'h0003,-16'h004e,-16'h000a,16'h003a,16'h0064,16'h0026,16'h0001,16'h0013,16'h0069,16'h003b,16'h0007,16'h0021,16'h0001,16'h0039,-16'h0008,16'h0039,16'h0022,-16'h0049,16'h0041,16'h0059,16'h0059,-16'h0045,-16'h0019,-16'h0012,16'h0029,-16'h0080,-16'h0080,-16'h0017,16'h0029,16'h0007,16'h0061,16'h002e,-16'h0015,-16'h000b,-16'h0019,16'h0031,16'h0054,16'h000f,16'h0011,16'h0002,-16'h00e2,16'h004c,-16'h003d,16'h000e,-16'h0019,16'h0002,16'h0025,16'h0075,-16'h0035,16'h004a,-16'h00a4,16'h0004,16'h008c,-16'h0011,-16'h00dd,16'h0014,-16'h0011,-16'h003a,-16'h000c,16'h0063,16'h0000,16'h000e,-16'h0097,16'h0087,16'h002b,-16'h0038,-16'h000c,16'h0035,16'h0049,16'h0002,16'h0015,16'h0010,16'h006e,16'h002f,-16'h000c,16'h0018,16'h0017,16'h002c,-16'h0005,16'h0057,16'h0011,-16'h0032,16'h003e,16'h006a,16'h0056,-16'h0023,-16'h0020,-16'h0034,16'h003a,-16'h0075,-16'h0077,16'h000a,16'h003d,16'h0002,16'h005f,16'h0059,16'h0004,-16'h0005,16'h0008,16'h001d,16'h0054,-16'h0004,-16'h0003,16'h0032,-16'h0104,16'h0030,-16'h003f,16'h0002,-16'h0016,-16'h0027,16'h0018,16'h0095,-16'h0022,16'h0036,-16'h0093,16'h0010,16'h00b6,16'h0038,-16'h00ad,16'h002c,16'h001b,-16'h001b,16'h000a,16'h0044,-16'h0001,16'h003c,-16'h0071,16'h007e,-16'h000e,-16'h001f,-16'h002f,16'h0048,16'h0003,-16'h0006,16'h0000,-16'h002c,16'h0083,16'h0028,-16'h001b,16'h004b,16'h0029,16'h0019,-16'h0004,16'h0068,16'h0024,-16'h0028,16'h0031,16'h0079,-16'h0010,-16'h0014,-16'h0056,-16'h003f,16'h004d,-16'h0066,-16'h007f,-16'h000a,16'h003e,16'h0010,16'h0048,16'h003d,16'h0006,16'h0004,16'h0003,16'h0008,16'h0065,16'h0005,-16'h0005,16'h004a,-16'h00e4,16'h0053,-16'h0019,-16'h0003,-16'h0003,-16'h0022,16'h0023,16'h0086,-16'h0026,16'h003e,-16'h0018,16'h0016,16'h009d,16'h0086,-16'h00a3,16'h0032,16'h0010,-16'h005c,16'h0015,16'h0062,16'h001e,16'h001f,-16'h004e,16'h0075,-16'h005d,-16'h0030,16'h000e,16'h0020,-16'h0022,-16'h000a,-16'h001d,-16'h0011,16'h0083,16'h003c,-16'h000d,16'h004c,16'h0041,16'h001c,-16'h001a,16'h0052,16'h0005,-16'h000e,16'h003d,16'h007a,-16'h0032,16'h001e,-16'h006d,-16'h003e,16'h0066,-16'h0062,-16'h005d,16'h0019,16'h0022,16'h0019,16'h0032,16'h0037,-16'h0009,-16'h0007,16'h0033,16'h0027,16'h0076,16'h0025,-16'h001c,16'h0060,-16'h0080,16'h0068,-16'h000c,16'h0019,16'h000f,16'h0009,16'h0022,16'h0086,-16'h0009,-16'h0009,16'h0018,16'h0018,16'h0097,16'h0093,-16'h009c,16'h0036,16'h0025,-16'h0098,16'h0021,16'h007d,16'h0059,16'h002a,16'h001e,16'h0007,-16'h005e,-16'h0017,16'h005e,16'h0008,-16'h000f,-16'h0011,-16'h0063,-16'h0016,16'h0064,16'h0048,-16'h0014,16'h0018,16'h003b,16'h001e,-16'h0017,16'h007a,-16'h001b,-16'h002b,16'h0028,16'h00a2,-16'h002f,16'h003b,-16'h003e,16'h0017,16'h0064,-16'h0058,-16'h006a,-16'h0017,16'h003d,-16'h000b,16'h001a,16'h0024,-16'h0022,-16'h0013,16'h001e,16'h001a,16'h004c,16'h0023,-16'h0017,16'h007a,-16'h001b,16'h005e,-16'h0005,16'h0043,-16'h0023,-16'h0020,16'h002f,16'h0097,16'h0023,-16'h0009,16'h005e,16'h0032,16'h0070,16'h0062,-16'h0081,16'h0026,16'h0022,-16'h00f4,16'h000b,16'h0034,16'h00a5,16'h003e,16'h000b,-16'h003d,-16'h0025,-16'h0028,16'h0078,16'h0016,-16'h0034,16'h0048,-16'h008a,-16'h0006,16'h005b,16'h004b,16'h003b,16'h0011,16'h0040,16'h003d,-16'h0050,16'h0089,16'h000c,-16'h000a,16'h0000,16'h007e,-16'h008b,16'h0047,-16'h003e,16'h002a,16'h0048,-16'h0009,-16'h0087,-16'h0034,16'h0047,-16'h0019,16'h0015,16'h0025,-16'h001b,16'h0000,16'h002f,16'h0017,16'h0034,16'h000e,-16'h001f,16'h0046,16'h002b,16'h003d,-16'h001b,16'h0075,-16'h001b,-16'h0007,16'h0049,16'h004c,16'h0032,-16'h0016,16'h007f,16'h0056,16'h0057,16'h0018,-16'h0068,16'h0022,16'h0041,-16'h00df,16'h0005,-16'h0066,16'h0080,16'h0034,16'h0022,-16'h0033,16'h0060,-16'h001d,-16'h000b,-16'h0008,-16'h002e,16'h0064,-16'h0058,-16'h0001,16'h0086,16'h0069,16'h0048,16'h003f,16'h0029,16'h0030,-16'h004e,16'h0099,16'h0011,16'h0005,-16'h0051,16'h0039,-16'h005a,16'h0028,-16'h0007,16'h000f,16'h0076,16'h0014,-16'h0062,-16'h0023,16'h003e,-16'h0010,16'h003a,16'h0038,16'h0019,16'h0008,16'h0017,16'h0031,16'h0043,16'h0013,-16'h0016,16'h0038,16'h0074,16'h0039,-16'h003c,16'h0066,-16'h001f,-16'h0010,16'h003e,16'h0027,16'h000f,-16'h0011,16'h0075,16'h0042,16'h0051,-16'h0084,-16'h0042,16'h0000,16'h0045,-16'h0001,16'h0035,-16'h009c,16'h005c,16'h0036,16'h0012,-16'h000f,16'h0052,16'h001d,-16'h009c,16'h000a,-16'h0021,16'h0076,-16'h0016,-16'h0004,16'h005a,16'h004c,16'h003d,16'h0012,16'h002d,16'h0009,-16'h0054,16'h0096,16'h001e,16'h0015,-16'h0040,16'h0003,16'h0025,16'h003c,16'h0027,-16'h000a,16'h0061,16'h000c,-16'h0070,-16'h0028,16'h0032,-16'h0006,16'h0021,16'h001c,16'h0037,16'h002a,-16'h0003,16'h003f,16'h0031,16'h001d,-16'h0028,16'h0027,16'h006f,16'h0049,-16'h0030,16'h0023,-16'h001c,-16'h002b,16'h0033,16'h0038,16'h0002,-16'h0019,16'h005e,-16'h001c,16'h0041,-16'h0086,-16'h0056,-16'h001e,16'h004b,16'h004b,16'h0046,-16'h0076,16'h002c,16'h0042,16'h000f,16'h0024,16'h0037,-16'h000f,-16'h00b5,-16'h0003,16'h0006,16'h0045,16'h0034,16'h0000,16'h0042,16'h004f,16'h0039,16'h001b,16'h0038,-16'h0006,-16'h0044,16'h0089,16'h004d,-16'h0038,-16'h0054,16'h000f,16'h004b,16'h0028,16'h001a,16'h001c,16'h0052,16'h000c,-16'h0072,-16'h004f,16'h0046,-16'h000d,16'h0024,16'h0032,16'h0033,16'h003c,-16'h0022,16'h0043,16'h0040,16'h000c,-16'h0035,16'h000a,16'h004a,16'h0030,-16'h000a,-16'h0004,-16'h000d,-16'h0002,16'h0048,16'h004b,-16'h000f,16'h0039,16'h001e,-16'h0043,16'h0065,-16'h0091,-16'h004f,-16'h002f,16'h005c,16'h0024,16'h0009,-16'h003b,-16'h002e,16'h002f,16'h003d,16'h0057,-16'h0008,16'h0018,-16'h0067,16'h000c,16'h0031,-16'h0002,16'h0004,16'h0026,16'h002a,16'h0030,16'h0039,16'h0020,16'h0019,16'h0007,-16'h0048,16'h0085,16'h0040,-16'h003a,-16'h0066,16'h0006,16'h008d,16'h0046,16'h002a,16'h001a,16'h0048,16'h0015,-16'h004a,-16'h0025,16'h005a,-16'h0014,16'h0034,16'h0028,16'h001e,16'h0024,-16'h0003,16'h001f,16'h003b,16'h0011,-16'h000f,-16'h0005,16'h004f,16'h002e,16'h001a,-16'h001e,-16'h0029,-16'h0020,16'h003f,16'h004f,16'h000b,16'h0024,-16'h0013,-16'h001e,16'h006e,-16'h006c,-16'h0055,16'h001e,16'h005e,16'h000c,-16'h0005,16'h0004,-16'h0076,16'h0036,16'h0027,16'h005b,-16'h001b,16'h0005,16'h0040,16'h000a,16'h000d,16'h002b,16'h0018,16'h001e,16'h0042,16'h004a,16'h0051,16'h000a,16'h0029,16'h001f,-16'h0025,16'h0061,16'h002c,-16'h0014,-16'h0038,-16'h0021,16'h007e,16'h0037,16'h006c,16'h0031,16'h0044,16'h0035,-16'h003d,-16'h0010,16'h0026,16'h0000,16'h0042,16'h002e,16'h0013,16'h0026,16'h0028,16'h0003,16'h000f,16'h000a,16'h0016,16'h0019,16'h0041,16'h0042,16'h0010,-16'h001d,-16'h0016,-16'h004e,16'h0035,16'h0042,16'h001d,16'h0015,-16'h0016,-16'h000d,16'h0078,-16'h0029,-16'h000d,16'h005f,16'h0061,-16'h000a,-16'h001a,16'h0012,-16'h0080,16'h001b,16'h003f,16'h0063,16'h0012,-16'h0007,16'h0060,16'h0001,16'h0002,16'h002e,16'h0020,16'h0031,16'h0032,16'h0040,16'h003a,16'h002a,16'h002a,16'h001e,-16'h0017,16'h0053,-16'h000d,-16'h0004,-16'h000b,-16'h000e,-16'h0029,16'h0022,16'h006f,16'h0021,16'h006a,16'h0054,-16'h0036,-16'h0019,16'h0022,16'h000b,16'h005e,16'h002b,16'h001b,16'h000e,16'h0017,16'h0001,-16'h0006,-16'h000c,-16'h0007,16'h0029,16'h0075,16'h0030,-16'h0015,16'h000a,-16'h0009,-16'h0063,16'h002b,16'h003b,16'h0016,16'h003d,-16'h0001,16'h0012,16'h0086,16'h0001,16'h000b,16'h006a,16'h005f,-16'h0044,-16'h0045,16'h002b,-16'h0065,16'h0028,16'h0045,16'h002e,16'h0025,16'h0003,16'h003a,16'h001f,-16'h0008,16'h0031,16'h001f,16'h002d,16'h0029,16'h003c,16'h0042,16'h0022,16'h001b,16'h001b,-16'h001e,16'h0061,-16'h0010,16'h0004,-16'h0015,-16'h0009,-16'h006e,16'h003c,16'h006e,16'h000b,16'h0064,16'h005e,-16'h0020,-16'h0001,16'h0017,16'h0023,16'h0069,16'h0016,16'h0028,16'h002d,-16'h0008,-16'h0010,-16'h0002,-16'h000b,-16'h0013,16'h0009,16'h0049,16'h0027,-16'h0008,-16'h0002,16'h0017,-16'h004a,16'h003f,16'h0031,16'h0028,16'h000b,-16'h001d,16'h0014,16'h005a,16'h0042,16'h000a,16'h007f,16'h004f,-16'h002e,-16'h0030,-16'h001b,-16'h0069,16'h000d,16'h001f,-16'h0014,16'h0030,16'h000a,16'h0022,16'h0012,-16'h0050,16'h0010,16'h0004,16'h0036,16'h001e,16'h0051,16'h000b,16'h0012,16'h0007,16'h0043,16'h000d,16'h006f,-16'h0008,16'h0015,16'h000f,-16'h0003,-16'h00aa,16'h0050,16'h006d,16'h0020,16'h0070,16'h004a,-16'h0010,-16'h0058,16'h003c,16'h0015,16'h005b,16'h003e,16'h001c,16'h001c,16'h001f,16'h0012,16'h000f,-16'h002e,16'h0017,16'h000d,16'h0025,16'h0039,-16'h0013,16'h0028,-16'h0008,-16'h0009,16'h005f,16'h004a,16'h0013,16'h0024,-16'h001d,16'h0021,16'h0010,16'h0049,-16'h001b,16'h0085,16'h0077,16'h0014,16'h0014,-16'h003a,-16'h004e,-16'h0018,-16'h000d,-16'h0009,16'h001d,16'h000d,-16'h000b,16'h0010,-16'h0044,16'h0031,16'h001b,16'h0042,16'h0025,16'h0022,-16'h0002,-16'h001e,-16'h0004,16'h003f,16'h002c,16'h006a,-16'h000e,16'h0017,-16'h0006,16'h0002,-16'h005d,16'h0038,16'h0064,16'h0024,16'h0068,16'h004b,-16'h000e,-16'h0072,16'h004d,-16'h0001,16'h005d,16'h001c,16'h0020,16'h0012,16'h0030,-16'h0003,16'h0013,-16'h002c,16'h0040,16'h0021,16'h000c,16'h0044,-16'h0011,16'h0012,16'h0000,-16'h0025,16'h006e,16'h0032,-16'h000c,16'h000f,-16'h0021,16'h0037,-16'h0004,16'h004d,-16'h000f,16'h006a,16'h0070,16'h0005,16'h002c,-16'h0053,-16'h0027,16'h0002,-16'h0017,-16'h0043,-16'h0004,16'h0024,16'h0005,-16'h000d,-16'h003a,16'h0026,16'h0044,16'h0031,16'h0058,16'h0011,16'h001f,-16'h001d,-16'h0006,16'h002e,16'h0025,16'h0082,-16'h002e,-16'h0005,16'h000a,16'h0018,-16'h0001,16'h0036,16'h0071,-16'h0005,16'h007c,16'h0033,-16'h000d,-16'h0054,16'h0046,16'h000c,16'h0060,16'h0009,16'h0033,16'h001c,16'h0038,-16'h0027,16'h0046,-16'h0032,16'h0013,16'h001b,16'h0003,16'h002b,-16'h000d,16'h0033,16'h0032,-16'h0019,16'h0062,16'h0023,-16'h0003,16'h0032,16'h0026,16'h002c,16'h0006,16'h004c,-16'h001f,16'h003d,16'h0076,-16'h001e,16'h0044,-16'h003d,16'h0001,16'h0023,16'h0006,-16'h0020,-16'h0022,16'h0009,-16'h0002,16'h0000,-16'h001e,16'h002b,16'h004e,16'h0032,16'h004e,16'h0028,16'h0038,16'h0002,16'h0035,16'h001a,-16'h0002,16'h007f,-16'h0029,-16'h0003,16'h001f,-16'h0020,16'h0023,16'h0045,16'h006c,-16'h001c,16'h006e,16'h001a,-16'h000d,-16'h0031,16'h0032,-16'h0001,16'h0030,-16'h0001,16'h001e,16'h0023,16'h0027,-16'h003b,16'h0038,-16'h0087,16'h0009,16'h0013,-16'h0004,16'h0035,-16'h001b,16'h002d,16'h003d,-16'h000d,16'h005c,16'h0024,-16'h0001,16'h0061,16'h0028,16'h0038,-16'h002e,16'h0046,-16'h0025,-16'h00d0,16'h006c,-16'h0020,16'h0081,-16'h001c,16'h002b,16'h002e,16'h0004,16'h002a,-16'h0032,16'h0010,-16'h0008,-16'h0026,-16'h0018,16'h001a,16'h004b,16'h001b,16'h003c,16'h0058,16'h0020,16'h0006,16'h0006,16'h001d,16'h0000,16'h005b,-16'h0016,-16'h0014,16'h0003,-16'h002e,16'h002c,16'h002c,16'h002d,-16'h003e,16'h007f,16'h0007,-16'h001b,16'h0000,16'h003f,-16'h0027,-16'h0027,16'h000d,16'h0016,16'h0031,16'h0013,-16'h004c,16'h0009,-16'h0105,-16'h0012,16'h0027,-16'h0041,16'h003e,-16'h0011,16'h0010,-16'h000c,16'h000c,16'h0052,16'h0021,16'h0030,16'h0057,16'h0033,16'h002e,-16'h0022,16'h0040,-16'h003e,-16'h0247,16'h005f,-16'h0023,16'h006c,16'h003a,16'h0037,16'h003f,-16'h0019,16'h0049,-16'h0041,16'h0012,-16'h001d,-16'h0030,16'h0016,16'h0053,16'h004b,16'h0054,16'h0033,16'h003c,-16'h001f,16'h0023,-16'h001c,16'h003b,16'h0015,16'h005e,-16'h000d,-16'h0022,-16'h0010,-16'h005f,16'h0000,16'h0032,16'h002f,-16'h0033,16'h0015,-16'h0022,16'h0010,16'h001a,16'h0042,-16'h0029,-16'h0020,-16'h000b,16'h0040,16'h0028,-16'h000b,-16'h0031,16'h001f,-16'h01b1,16'h001a,16'h001d,16'h0005,16'h0036,16'h000d,-16'h0015,16'h001c,-16'h0006,16'h003a,-16'h0001,16'h001a,-16'h004b,16'h0029,-16'h0029,-16'h0029,16'h001e,-16'h007c,-16'h029b,16'h004a,-16'h0005,16'h0075,16'h0010,16'h0032,16'h0020,-16'h000a,16'h005d,-16'h003e,-16'h000e,16'h0011,-16'h0020,16'h0028,16'h0043,16'h0054,16'h0041,16'h0031,16'h0032,-16'h0031,-16'h0003,-16'h0006,16'h001d,-16'h0016,16'h0074,-16'h001f,-16'h003a,-16'h001a,-16'h0063,16'h0003,16'h0024,16'h0012,-16'h000b,-16'h0113,-16'h001c,16'h0001,-16'h0006,16'h0029,-16'h002d,16'h000e,-16'h0018,16'h001a,16'h0047,-16'h002f,-16'h003f,16'h001b,-16'h01c1,16'h0018,16'h002f,16'h0022,16'h0005,16'h0033,-16'h000f,16'h0008,-16'h003b,16'h0054,-16'h0007,-16'h0006,-16'h00be,16'h0032,-16'h008f,-16'h0043,-16'h004b,-16'h0038,-16'h016f,16'h004b,-16'h0007,16'h005e,-16'h003d,16'h002a,16'h001f,-16'h002c,16'h006a,-16'h0026,-16'h0036,16'h002e,-16'h001a,16'h0025,16'h0035,16'h0011,16'h0058,16'h0052,16'h0012,-16'h003e,16'h0039,16'h0012,16'h001a,-16'h0004,16'h0044,-16'h0018,16'h000c,-16'h0032,-16'h001b,16'h003b,16'h003e,16'h0012,16'h0006,-16'h022f,16'h0025,-16'h000b,-16'h002b,16'h000d,-16'h0045,16'h002a,-16'h0027,16'h001e,16'h003c,-16'h003a,-16'h0046,16'h0061,-16'h0178,16'h0049,16'h0075,16'h0059,16'h002c,16'h002b,-16'h0021,-16'h002e,-16'h0044,16'h0038,16'h0011,16'h0003,-16'h0097,-16'h000e,-16'h00d6,-16'h005e,-16'h004f,-16'h0023,-16'h00ca,16'h003c,16'h0002,-16'h00d3,-16'h003c,-16'h000c,16'h0006,-16'h0057,16'h0074,16'h0016,-16'h000b,16'h004a,-16'h003e,16'h0026,-16'h000d,16'h0001,16'h0068,16'h0058,16'h002d,-16'h0078,16'h0040,16'h0008,16'h0016,16'h002c,16'h001e,16'h0000,16'h000f,-16'h0004,-16'h0007,16'h001f,16'h0011,16'h0010,16'h003b,-16'h01a6,16'h003c,-16'h0024,-16'h0036,16'h0012,-16'h0031,16'h0049,-16'h0038,16'h0019,-16'h0007,-16'h002b,-16'h003a,-16'h0001,-16'h00fd,16'h0058,16'h00a9,16'h0061,16'h0013,16'h0032,-16'h0030,-16'h0025,-16'h0019,16'h005a,16'h0016,-16'h0018,-16'h0081,-16'h002c,-16'h00e0,-16'h0037,-16'h001a,-16'h0046,-16'h0065,16'h0056,-16'h0016,-16'h01c8,-16'h0026,-16'h0066,16'h0025,-16'h003f,16'h0034,16'h0038,16'h0000,16'h0029,-16'h0032,16'h0025,16'h000b,-16'h0002,16'h009b,16'h0058,16'h001f,-16'h00a0,16'h0014,-16'h0015,-16'h0009,16'h0048,16'h0017,16'h0006,-16'h0004,16'h0026,-16'h0003,16'h000c,-16'h0006,16'h001f,16'h002a,-16'h00cf,16'h0020,16'h000e,-16'h0056,16'h0037,-16'h001b,16'h0049,-16'h0013,16'h0039,-16'h0083,16'h0005,-16'h0041,-16'h0056,-16'h00d7,16'h003f,16'h0092,16'h003e,16'h000c,16'h0031,16'h0000,-16'h0035,16'h0007,16'h0054,16'h0009,16'h0020,-16'h003b,-16'h0056,-16'h00ae,-16'h0056,-16'h0009,-16'h0022,-16'h0018,16'h003f,-16'h0002,-16'h018f,-16'h0006,-16'h0085,-16'h0009,-16'h0011,16'h003a,16'h001c,16'h002c,16'h0005,16'h0000,16'h0012,16'h000d,-16'h0006,16'h0089,16'h005f,16'h000c,-16'h009c,-16'h000e,-16'h001c,16'h000f,16'h007b,16'h0009,16'h0037,16'h000d,16'h0049,16'h0025,16'h000c,16'h0016,16'h0022,16'h0025,-16'h004f,-16'h0027,-16'h0001,-16'h0011,16'h003d,16'h0003,16'h003e,-16'h001f,16'h002c,-16'h0095,-16'h0025,-16'h003e,-16'h0037,-16'h00b8,16'h0000,16'h0053,16'h0042,16'h000a,16'h0060,16'h0028,-16'h0046,16'h000b,16'h0045,16'h0013,16'h001a,-16'h001b,-16'h0076,-16'h0075,-16'h0049,16'h0008,-16'h0050,16'h0030,16'h0077,16'h0010,-16'h0115,-16'h0015,-16'h00b5,16'h004b,-16'h0022,16'h001b,16'h000a,16'h0047,16'h0013,16'h0024,16'h0006,16'h0004,16'h0028,16'h0068,16'h00a4,-16'h0024,-16'h0096,-16'h000a,-16'h001a,-16'h0015,16'h0036,16'h0033,16'h001f,16'h0017,16'h0070,16'h0007,16'h0000,16'h0023,16'h0023,16'h0039,-16'h0020,-16'h0094,-16'h0027,16'h001d,16'h005c,16'h0022,16'h005e,16'h0049,-16'h0017,-16'h0014,16'h003f,16'h0043,16'h0042,16'h0051,-16'h0013,16'h00f1,-16'h0042,16'h0082,16'h0019,16'h0008,16'h0015,16'h0000,-16'h001e,16'h0020,-16'h002f,-16'h004a,16'h0008,16'h0099,16'h0009,-16'h0014,-16'h0082,-16'h0032,-16'h002c,-16'h003e,16'h001c,16'h00e3,16'h007e,16'h0037,16'h002c,-16'h005b,-16'h001d,16'h0039,-16'h0015,-16'h0015,16'h009f,-16'h0009,16'h0025,16'h005c,16'h0017,-16'h0006,-16'h000e,16'h001c,-16'h0004,16'h0049,-16'h003c,16'h003d,-16'h0023,-16'h0015,16'h0021,-16'h004b,16'h002a,16'h0017,-16'h0049,-16'h001d,-16'h0022,-16'h0003,-16'h0029,16'h0052,16'h0021,16'h0010,16'h0058,16'h007b,-16'h0021,-16'h0034,16'h0021,16'h004c,16'h0012,16'h0050,16'h002c,16'h00a8,-16'h005b,16'h0083,16'h001a,16'h0013,16'h0019,16'h0026,-16'h002b,16'h0013,-16'h003f,-16'h0025,16'h0012,16'h0003,16'h002a,-16'h001b,-16'h00bc,-16'h002e,-16'h002f,-16'h0029,-16'h0018,16'h00bf,16'h0091,16'h0048,16'h0042,-16'h0077,-16'h002a,-16'h000e,-16'h001f,16'h002a,16'h00a7,-16'h0002,16'h0013,16'h0023,16'h004a,-16'h0003,-16'h000d,16'h001c,-16'h002e,16'h002e,-16'h0037,16'h0016,-16'h0029,-16'h0023,16'h0031,16'h0000,16'h0071,-16'h0008,-16'h0017,16'h0009,-16'h001c,-16'h0002,-16'h0017,16'h0022,16'h002e,16'h0025,16'h0058,16'h0075,-16'h0055,-16'h001c,16'h000c,16'h000e,-16'h001e,16'h0043,16'h0042,16'h007e,-16'h006c,16'h004b,16'h0013,16'h0027,-16'h0003,16'h0039,16'h0003,16'h0024,-16'h0028,-16'h001c,-16'h001d,-16'h0003,16'h0071,-16'h001b,-16'h0110,-16'h000b,-16'h001c,-16'h0051,-16'h0028,16'h0076,16'h0046,16'h0029,16'h0017,-16'h001b,16'h0001,-16'h0051,-16'h0011,16'h0018,16'h007d,-16'h0001,-16'h0019,16'h0033,16'h0051,16'h001e,-16'h000b,16'h0020,-16'h0032,16'h000f,-16'h0048,16'h001e,16'h0012,-16'h0039,16'h0032,16'h001c,16'h0080,-16'h0018,-16'h0034,-16'h003d,-16'h0011,16'h0001,-16'h0042,16'h001d,16'h004a,16'h0026,16'h0063,16'h004e,-16'h0087,16'h0007,16'h0011,16'h0006,-16'h0018,16'h0011,16'h002e,16'h0033,-16'h009e,16'h002a,-16'h0047,16'h0017,-16'h000f,16'h0003,-16'h0007,16'h002e,-16'h002f,16'h0015,-16'h006d,-16'h0015,16'h0086,-16'h000f,-16'h00fa,16'h0009,-16'h0028,-16'h002e,-16'h002b,16'h0078,-16'h0017,16'h0028,-16'h0022,16'h002a,16'h0017,-16'h0043,-16'h002f,16'h002c,16'h0044,16'h000f,-16'h0017,16'h0048,16'h006b,16'h0011,-16'h0003,16'h0022,16'h000b,16'h001e,-16'h001b,16'h0036,16'h000a,-16'h0033,16'h0063,16'h008c,16'h0062,-16'h002a,-16'h0037,-16'h002f,16'h001b,-16'h0001,-16'h0052,16'h001a,16'h0034,16'h0023,16'h0070,16'h002c,-16'h0071,16'h000c,-16'h000a,16'h001a,16'h0002,-16'h0006,16'h002f,16'h002b,-16'h00b4,16'h0006,-16'h002a,16'h0003,16'h000b,-16'h0005,16'h0017,16'h004d,-16'h0038,16'h0026,-16'h00a1,-16'h000e,16'h007b,16'h0014,-16'h0092,16'h001e,-16'h0028,16'h0000,-16'h0016,16'h0064,16'h0003,16'h0014,-16'h008c,16'h0073,16'h001e,-16'h0058,-16'h0024,16'h0041,16'h0051,-16'h0012,16'h000c,16'h0019,16'h008b,16'h0010,16'h001c,16'h002b,16'h0037,16'h002a,-16'h0004,16'h005a,16'h001a,-16'h0012,16'h0024,16'h0088,16'h0019,-16'h0031,-16'h004f,-16'h0035,16'h0016,16'h0020,-16'h007a,16'h0018,16'h0033,16'h000a,16'h004b,16'h005f,-16'h007b,16'h0037,16'h0006,16'h0009,16'h001d,-16'h0004,16'h003a,16'h003f,-16'h00a6,16'h0029,-16'h000a,-16'h0023,-16'h000e,-16'h001e,16'h0002,16'h0045,-16'h0032,16'h0037,-16'h008a,16'h0024,16'h008c,16'h005e,-16'h0059,16'h0041,-16'h0012,-16'h0015,-16'h0003,16'h0078,-16'h0001,16'h0025,-16'h0080,16'h0072,-16'h0028,-16'h0069,-16'h003f,16'h0013,16'h003d,-16'h0038,16'h001a,-16'h0011,16'h0084,16'h001c,16'h0000,16'h003a,16'h0028,16'h000d,-16'h0026,16'h0062,16'h0036,16'h0006,16'h0028,16'h0084,-16'h0017,-16'h001a,-16'h0046,-16'h0040,16'h004b,16'h000c,-16'h007e,16'h001a,16'h004e,16'h0017,16'h0054,16'h0038,-16'h005c,16'h0027,16'h001b,16'h0026,16'h0060,-16'h0016,16'h0014,16'h0045,-16'h009a,16'h004c,16'h0012,-16'h0014,-16'h0004,-16'h0025,16'h0021,16'h006c,-16'h0016,16'h0033,-16'h0031,16'h0023,16'h00b4,16'h007b,-16'h007d,16'h003d,-16'h0010,-16'h0023,16'h0021,16'h0060,16'h0016,16'h0038,-16'h002b,16'h0049,-16'h0066,-16'h0032,16'h0005,16'h000d,-16'h002f,-16'h0003,-16'h000b,-16'h0022,16'h0064,16'h0009,-16'h0026,16'h002c,16'h0011,16'h001b,-16'h0036,16'h005c,16'h0022,16'h0016,16'h002a,16'h0095,-16'h004d,-16'h000c,-16'h0061,-16'h0032,16'h000d,16'h0031,-16'h0067,16'h002c,16'h0017,16'h0015,16'h0053,16'h0052,-16'h00a7,16'h000d,16'h000e,16'h0007,16'h0058,-16'h0005,16'h001f,16'h0043,-16'h003c,16'h0040,-16'h0007,16'h001c,16'h0014,-16'h0032,16'h0031,16'h003f,-16'h002b,16'h000d,16'h000c,16'h002d,16'h0093,16'h0064,-16'h0070,16'h0027,-16'h0006,-16'h0093,16'h0023,16'h009c,16'h007c,16'h0052,16'h001c,-16'h0003,-16'h0057,-16'h003d,16'h0034,-16'h0002,-16'h0055,16'h0011,-16'h0062,-16'h0004,16'h003a,-16'h0001,-16'h0019,16'h0034,16'h001a,16'h0037,-16'h005d,16'h0065,16'h0000,16'h0028,16'h0016,16'h0090,-16'h007f,16'h000e,-16'h006f,-16'h0007,16'h002c,16'h0051,-16'h006f,-16'h0002,16'h0029,16'h0005,16'h0040,16'h0056,-16'h0096,-16'h0008,16'h0056,16'h0027,16'h002b,16'h0011,16'h0025,16'h004b,16'h0011,16'h005b,-16'h0009,16'h0043,-16'h000a,-16'h002e,16'h0030,16'h003c,16'h0013,-16'h0033,16'h0047,16'h0039,16'h008a,16'h003f,-16'h0055,16'h0016,-16'h0007,-16'h00a7,-16'h0009,16'h004f,16'h0073,16'h003f,16'h000e,-16'h0045,-16'h0015,-16'h002a,16'h0053,16'h000c,-16'h002c,16'h006f,-16'h0069,-16'h0022,16'h0067,16'h003b,16'h0004,16'h0026,16'h003c,16'h0016,-16'h0051,16'h0050,-16'h0006,16'h0032,-16'h0018,16'h0081,-16'h007f,16'h0020,-16'h0069,16'h000a,16'h0011,16'h0061,-16'h0084,-16'h000a,16'h0026,-16'h0006,16'h004e,16'h0026,-16'h0071,-16'h0001,16'h0055,16'h003d,16'h0017,16'h001e,-16'h000b,16'h0050,16'h002f,16'h006e,-16'h0038,16'h0038,-16'h0007,-16'h0047,16'h0038,16'h0030,16'h001e,-16'h0024,16'h0052,16'h0057,16'h0086,-16'h003b,-16'h004d,16'h001e,16'h0017,-16'h004c,16'h0029,-16'h0034,16'h005b,16'h0030,16'h001a,-16'h001d,16'h004f,-16'h000e,-16'h0058,16'h0001,-16'h0008,16'h0054,-16'h005d,-16'h0035,16'h0070,16'h0030,16'h0044,16'h0026,16'h002d,16'h001a,-16'h003c,16'h005b,-16'h0013,16'h0046,-16'h005e,16'h004d,-16'h003f,16'h001f,-16'h0028,16'h000e,16'h002f,16'h007b,-16'h006f,-16'h002c,16'h0031,-16'h000e,16'h005f,16'h003c,-16'h0044,16'h002f,16'h0036,16'h0026,-16'h0004,16'h0018,16'h000f,16'h0040,16'h004a,16'h0045,-16'h002c,16'h0051,-16'h0023,-16'h0032,16'h004a,16'h000c,16'h0024,-16'h0021,16'h006c,16'h0020,16'h0049,-16'h0090,-16'h0065,16'h000b,16'h0020,16'h002f,16'h002e,-16'h008f,16'h0027,16'h0044,16'h0030,-16'h001e,16'h003c,-16'h0004,-16'h00c3,-16'h0005,-16'h0020,16'h003e,-16'h0017,-16'h0039,16'h0059,16'h0046,16'h004d,16'h0020,16'h002e,-16'h0010,-16'h001f,16'h0072,16'h0025,16'h0032,-16'h002e,16'h002a,16'h0026,16'h0013,16'h0015,16'h0010,16'h0031,16'h0057,-16'h0059,-16'h0029,16'h0045,-16'h000b,16'h003f,16'h004e,-16'h0029,16'h0024,16'h0049,16'h0036,16'h000a,16'h0025,16'h000a,16'h001f,16'h0057,16'h0048,-16'h0026,16'h0017,-16'h0020,-16'h0029,16'h0050,16'h0014,16'h0009,-16'h0006,16'h0043,-16'h0029,16'h005e,-16'h00a2,-16'h0067,16'h0005,16'h0015,16'h0078,16'h0029,-16'h00ad,-16'h001c,16'h0052,16'h000a,16'h0045,16'h0014,-16'h0009,-16'h00ba,16'h0004,-16'h0008,16'h0015,-16'h0003,-16'h000a,16'h0053,16'h0038,16'h003a,16'h0029,16'h0046,16'h0004,-16'h002c,16'h008f,16'h0019,-16'h0011,-16'h005b,16'h000c,16'h006e,16'h000c,16'h000d,16'h0040,16'h000b,16'h0043,-16'h0060,-16'h0067,16'h0034,16'h0000,16'h0031,16'h0033,-16'h004d,16'h0014,16'h0020,16'h0010,16'h0036,16'h000d,16'h0014,16'h0017,16'h0039,16'h0052,-16'h0013,-16'h0009,-16'h002d,-16'h0002,16'h0045,16'h001d,16'h0002,16'h0049,-16'h0002,-16'h0024,16'h0079,-16'h006c,-16'h005e,-16'h000b,16'h0035,16'h003c,-16'h0002,-16'h0093,-16'h007d,16'h0038,16'h0010,16'h0062,16'h000c,16'h0002,-16'h0056,-16'h0026,16'h0008,16'h0024,16'h001e,16'h000f,16'h0025,16'h002f,16'h003f,16'h002f,16'h0027,-16'h0015,-16'h003f,16'h0081,16'h003b,-16'h0003,-16'h005b,-16'h0003,16'h009b,16'h0006,16'h0007,16'h003a,16'h000e,16'h001f,-16'h0060,-16'h005a,16'h004f,16'h0002,16'h002b,16'h0040,-16'h0046,16'h001c,16'h0035,-16'h0011,16'h002a,16'h000d,16'h001e,16'h001c,16'h0035,16'h0053,16'h0009,-16'h0016,-16'h001a,-16'h0010,16'h0046,16'h0034,16'h000a,16'h0049,-16'h0026,-16'h002c,16'h0060,-16'h004a,-16'h0064,16'h001b,16'h003d,16'h0038,-16'h000a,-16'h005d,-16'h0077,16'h003f,16'h0038,16'h004c,16'h001b,16'h0019,16'h003e,-16'h0034,16'h0017,16'h0020,16'h0002,16'h002c,16'h001b,16'h0062,16'h0058,16'h003a,16'h002e,-16'h0008,-16'h003f,16'h0077,16'h002c,16'h0013,-16'h0057,-16'h0001,16'h0062,16'h0003,16'h0045,16'h0033,16'h0015,16'h002c,-16'h0080,-16'h0049,16'h001b,16'h0009,16'h0044,16'h0042,-16'h0036,16'h000f,16'h001c,-16'h0015,16'h0010,16'h0000,16'h0017,16'h002f,16'h004c,16'h004d,-16'h0002,-16'h0027,-16'h0002,-16'h0021,16'h002e,16'h003e,16'h0039,16'h003e,-16'h001e,-16'h0004,16'h006d,16'h0018,-16'h0040,16'h0052,16'h0060,16'h000d,16'h0005,-16'h000f,-16'h006e,16'h003b,16'h0058,16'h0000,16'h0042,-16'h000d,16'h0061,-16'h0027,16'h0005,16'h0023,16'h0005,16'h002b,16'h000c,16'h0046,16'h003c,16'h0048,16'h0012,16'h0015,-16'h0019,16'h0076,16'h001b,-16'h0015,-16'h0027,-16'h0034,-16'h0026,-16'h0011,16'h006f,16'h0039,16'h0029,16'h0033,-16'h0061,-16'h004c,16'h0020,16'h0004,16'h005a,16'h0030,-16'h003b,16'h0033,16'h000b,-16'h0036,-16'h0001,-16'h000e,16'h0002,16'h0034,16'h0043,16'h0070,-16'h001d,-16'h0012,-16'h000e,-16'h003b,16'h002c,16'h0039,16'h0028,16'h0043,-16'h0004,-16'h000c,16'h0078,16'h003c,16'h000b,16'h0066,16'h007b,-16'h003c,-16'h0016,-16'h0005,-16'h0046,16'h0035,16'h005e,-16'h0001,16'h0015,-16'h0013,16'h002c,-16'h0001,16'h000d,16'h002d,16'h0000,16'h0045,16'h0007,16'h004c,16'h0036,16'h0014,16'h0027,16'h0042,-16'h0023,16'h0072,16'h0015,16'h0044,-16'h000c,-16'h0033,-16'h0081,16'h0000,16'h0048,16'h0027,16'h0017,16'h003c,-16'h0054,-16'h0033,16'h002f,16'h0035,16'h0085,16'h0045,-16'h0062,16'h0020,16'h001a,-16'h002f,-16'h0021,-16'h005b,16'h0002,16'h002c,16'h0029,16'h005c,-16'h0009,16'h0005,16'h0001,-16'h0018,16'h004b,16'h001f,16'h001c,16'h0033,-16'h002c,16'h0009,16'h003a,16'h0026,16'h0000,16'h0096,16'h0062,-16'h0039,-16'h000f,-16'h002d,-16'h0028,16'h0010,16'h0028,-16'h002c,16'h002d,-16'h0017,16'h0020,-16'h0008,16'h0001,16'h0040,-16'h0011,16'h0033,-16'h0007,16'h0016,16'h0000,16'h0012,16'h0019,16'h003f,-16'h0008,16'h008c,-16'h000d,16'h004b,16'h001e,-16'h002f,-16'h00b6,16'h0031,16'h0025,16'h000b,16'h004e,16'h0049,-16'h0059,-16'h0031,16'h0054,16'h0028,16'h0087,16'h0038,-16'h0029,16'h0014,16'h0004,-16'h003f,16'h000b,-16'h0053,-16'h0004,16'h001e,16'h0010,16'h0048,-16'h0023,16'h000f,-16'h0013,-16'h0005,16'h0057,16'h0018,16'h001c,16'h002f,-16'h0034,16'h0024,16'h0016,16'h005c,-16'h0027,16'h0096,16'h0073,16'h0000,16'h001f,-16'h0050,-16'h000c,16'h0030,16'h001a,-16'h0035,-16'h0008,-16'h0011,-16'h0001,-16'h000e,16'h000e,16'h0032,16'h001a,16'h0025,16'h0008,16'h0021,16'h000e,16'h0003,-16'h000d,16'h0031,-16'h000a,16'h007b,-16'h0013,16'h0040,16'h0001,-16'h002e,-16'h0065,16'h0011,16'h003c,16'h0016,16'h0046,16'h004f,-16'h0069,-16'h0051,16'h0050,16'h0005,16'h0066,16'h003f,-16'h002e,16'h001c,16'h0039,-16'h0065,16'h0024,-16'h0081,16'h0000,16'h001c,16'h001c,16'h0065,-16'h000d,-16'h0004,-16'h0006,16'h0008,16'h005a,16'h0027,16'h0002,16'h0024,-16'h0004,16'h0057,16'h0037,16'h003a,-16'h0009,16'h0084,16'h0081,16'h0001,16'h0050,-16'h0032,-16'h0001,16'h0022,16'h000f,-16'h000f,-16'h0037,16'h0000,-16'h0029,16'h0008,-16'h001a,16'h001a,16'h005d,16'h0041,16'h0014,-16'h000a,-16'h0005,16'h0031,16'h000f,16'h004a,16'h0026,16'h0057,-16'h0011,16'h0023,16'h0012,-16'h0039,16'h0005,16'h0006,16'h0043,-16'h001a,16'h0056,16'h0052,-16'h0092,-16'h0031,16'h0056,16'h0012,16'h0074,16'h001c,-16'h0014,16'h0002,16'h0033,-16'h0059,16'h003f,-16'h00e4,-16'h000b,16'h0030,16'h000a,16'h0061,-16'h0010,16'h001d,-16'h0007,16'h0002,16'h0050,16'h0009,16'h0001,16'h001a,16'h002a,16'h002c,16'h0034,16'h0034,-16'h0023,16'h0043,16'h006b,-16'h000b,16'h0057,-16'h0031,16'h001d,16'h002f,-16'h0018,16'h0000,-16'h0038,16'h0010,-16'h000d,-16'h0018,-16'h003d,16'h0044,16'h003a,16'h0038,16'h0039,16'h0010,16'h000e,16'h0033,16'h0000,16'h004b,16'h000b,16'h0047,-16'h0012,16'h0005,16'h0027,-16'h0031,16'h002d,16'h0020,16'h0040,-16'h001a,16'h0053,16'h0024,-16'h00a5,16'h000a,16'h0017,16'h0023,16'h003e,16'h0015,16'h0004,16'h004a,16'h0005,-16'h0053,16'h0017,-16'h016c,-16'h000c,16'h0032,-16'h000b,16'h003b,16'h000a,16'h003f,16'h001b,16'h0018,16'h0044,16'h0030,-16'h0006,16'h0065,16'h0023,16'h0013,16'h001a,16'h002d,-16'h0005,-16'h00ad,16'h0077,-16'h0005,16'h0068,-16'h001d,16'h0030,16'h0056,-16'h0015,16'h0021,-16'h0031,16'h000f,-16'h0011,-16'h0021,16'h0000,16'h001e,16'h001a,16'h003d,16'h0046,16'h0032,-16'h0041,16'h003e,-16'h000e,16'h002a,-16'h0008,16'h003a,16'h000b,16'h0001,16'h0001,-16'h0034,16'h0038,16'h0026,16'h001e,-16'h0034,16'h0042,16'h001b,-16'h0072,16'h0028,-16'h000b,16'h0001,16'h0000,-16'h000b,16'h0025,16'h005d,-16'h0012,-16'h0038,16'h0018,-16'h01c6,-16'h000e,16'h0033,-16'h0008,16'h0037,16'h0007,16'h002a,16'h0030,16'h0016,16'h0029,16'h0035,16'h0007,16'h0034,16'h0039,-16'h001e,16'h000c,16'h001e,-16'h0039,-16'h025d,16'h0041,16'h0001,16'h0069,16'h0000,16'h0022,16'h005e,-16'h001f,16'h006a,-16'h0033,16'h0009,-16'h001e,-16'h0046,16'h0009,16'h0013,16'h0011,16'h003f,16'h002f,16'h0043,-16'h005f,16'h0029,-16'h0033,16'h0033,-16'h0027,16'h0083,16'h0015,-16'h001c,-16'h000c,-16'h003b,16'h0009,16'h0021,16'h0034,-16'h0041,-16'h0016,-16'h0006,-16'h0052,16'h0008,16'h0020,-16'h000f,-16'h0007,-16'h0019,16'h000f,16'h0059,-16'h001a,-16'h0027,16'h002b,-16'h01b2,16'h0022,16'h0031,-16'h0005,16'h0020,16'h001e,16'h0003,16'h000d,-16'h0025,16'h0032,16'h0016,16'h002c,-16'h0078,16'h0011,-16'h006e,16'h000e,-16'h0031,-16'h0070,-16'h02b8,16'h0056,-16'h000c,16'h007e,-16'h000f,16'h0018,16'h0040,16'h0016,16'h0060,-16'h0020,-16'h0002,16'h0013,-16'h004f,16'h0000,16'h0020,16'h0015,16'h005e,16'h0030,16'h0025,-16'h0099,16'h0025,-16'h0008,16'h0039,-16'h000f,16'h006b,-16'h000a,-16'h0008,-16'h0025,-16'h0035,-16'h0010,16'h001b,16'h002b,-16'h0020,-16'h0199,-16'h000e,-16'h005e,-16'h0024,16'h0027,-16'h003e,16'h002a,16'h0014,16'h001e,16'h005c,-16'h0039,-16'h0038,16'h003e,-16'h015c,16'h0032,16'h0039,16'h0000,16'h0004,16'h002d,-16'h002d,-16'h0002,-16'h0045,16'h0032,16'h0013,16'h0008,-16'h00ce,16'h0006,-16'h00cc,16'h0005,-16'h0066,-16'h002a,-16'h0172,16'h0062,16'h0001,16'h0055,-16'h005d,-16'h0014,16'h0026,16'h000b,16'h0070,16'h0000,-16'h0025,16'h004e,-16'h001d,16'h001c,16'h0009,16'h000a,16'h0043,16'h0009,16'h0013,-16'h008f,16'h002d,16'h000a,16'h0010,16'h000d,16'h005d,-16'h0011,16'h001c,-16'h0016,-16'h000d,16'h0006,16'h0016,16'h0047,-16'h000b,-16'h0276,-16'h0001,-16'h0039,-16'h001b,16'h0000,-16'h0051,16'h0043,16'h0011,16'h001e,16'h0040,-16'h0035,-16'h0029,16'h0038,-16'h00f0,16'h001c,16'h0072,16'h0040,16'h0005,16'h0039,-16'h0041,-16'h0033,-16'h002a,16'h0027,16'h0020,-16'h0018,-16'h008b,-16'h000b,-16'h0104,-16'h0010,-16'h0078,-16'h0027,-16'h00b7,16'h0049,-16'h0007,-16'h00d1,-16'h0064,-16'h0054,16'h0033,-16'h001d,16'h0071,-16'h0001,-16'h0028,16'h004b,-16'h004a,16'h0023,16'h0006,-16'h001f,16'h0071,16'h0045,-16'h0005,-16'h00db,16'h002c,-16'h0018,16'h0018,16'h0037,16'h0037,16'h000e,16'h000a,16'h001f,-16'h000f,16'h003b,16'h0008,16'h0015,16'h002f,-16'h018e,16'h0045,-16'h005c,-16'h0027,16'h003e,-16'h002b,16'h0067,-16'h0005,16'h0022,16'h0025,-16'h001b,-16'h0030,-16'h0005,-16'h00c2,16'h002a,16'h00a5,16'h0043,-16'h0016,16'h003a,-16'h000d,-16'h0034,16'h000d,16'h0051,-16'h0005,-16'h0001,-16'h007a,-16'h0028,-16'h00c5,-16'h0007,-16'h001d,-16'h0026,-16'h005d,16'h007c,16'h001a,-16'h01b8,-16'h002e,-16'h009a,16'h001a,-16'h0017,16'h0059,16'h0010,-16'h0004,16'h002a,-16'h0038,16'h0003,16'h0011,-16'h0016,16'h008f,16'h0018,16'h0013,-16'h00e8,16'h0007,-16'h0013,-16'h0005,16'h006f,16'h0019,16'h0041,16'h002d,16'h0046,-16'h0005,16'h002c,-16'h000f,16'h0017,16'h0014,-16'h00c2,16'h0033,-16'h004d,-16'h001e,16'h0043,-16'h0025,16'h006b,16'h0017,16'h0014,-16'h0053,-16'h002d,-16'h002c,-16'h0055,-16'h00cd,16'h0007,16'h00a5,16'h0023,-16'h0028,16'h005c,16'h0010,-16'h0055,16'h0015,16'h002c,-16'h0006,16'h0002,-16'h003e,-16'h002a,-16'h0097,-16'h0012,-16'h0028,-16'h0019,-16'h0013,16'h0065,-16'h000a,-16'h0182,-16'h000b,-16'h008b,16'h0000,-16'h001f,16'h0052,16'h0027,16'h0024,16'h000a,-16'h0011,16'h0011,16'h0003,-16'h0017,16'h0070,16'h0044,-16'h0002,-16'h0087,-16'h002c,-16'h0027,-16'h0010,16'h0084,16'h003d,16'h0058,16'h0033,16'h006c,16'h0020,16'h0023,-16'h0018,16'h001f,16'h002d,-16'h003d,-16'h001f,-16'h0046,16'h0013,16'h0007,-16'h002a,16'h004c,16'h0029,16'h0010,-16'h00ab,-16'h003f,-16'h005a,-16'h0063,-16'h009b,16'h0007,16'h008f,16'h0044,16'h0013,16'h0039,16'h0031,-16'h006c,16'h0028,16'h0063,16'h0015,16'h001e,-16'h0046,-16'h003e,-16'h0071,-16'h000c,-16'h0028,-16'h0041,16'h0038,16'h0078,16'h0033,-16'h011a,-16'h000c,-16'h009a,16'h0030,-16'h0033,16'h0000,16'h001e,16'h0065,16'h0008,16'h0030,16'h0031,-16'h0013,16'h004e,16'h004e,16'h0069,-16'h0012,-16'h008d,-16'h0008,-16'h0019,-16'h001a,16'h005d,16'h0047,16'h0016,16'h000f,16'h006e,16'h0012,-16'h0007,-16'h0017,16'h0002,16'h0012,16'h0000,-16'h0043,-16'h0039,16'h0021,16'h0062,16'h0044,16'h004d,16'h0020,-16'h004d,16'h0007,16'h003f,16'h0021,16'h004f,16'h0074,-16'h003b,16'h00ae,-16'h003a,16'h0099,16'h0015,-16'h0004,16'h000b,16'h000e,-16'h0010,16'h002b,-16'h005a,-16'h0019,16'h0017,16'h00a6,-16'h0007,-16'h0020,-16'h0098,-16'h0014,-16'h0004,-16'h0002,-16'h000c,16'h00f1,16'h0073,16'h0050,16'h0037,-16'h0068,-16'h002f,16'h0040,-16'h0018,-16'h0002,16'h00a5,-16'h000e,16'h0007,16'h0044,16'h000a,-16'h0007,-16'h0003,16'h000d,16'h0028,16'h0038,-16'h0025,16'h005b,-16'h0026,-16'h000d,16'h0028,-16'h0041,16'h003e,16'h000d,-16'h0042,-16'h0044,-16'h003b,16'h0045,-16'h001a,16'h0058,16'h005e,16'h0026,16'h002e,16'h006e,-16'h0046,-16'h0022,16'h002b,16'h0012,16'h0033,16'h004c,16'h0022,16'h00b6,-16'h0083,16'h006f,16'h000c,-16'h000d,16'h0006,16'h0036,-16'h0023,16'h0042,-16'h003c,-16'h0030,16'h0019,16'h0029,16'h0014,-16'h000a,-16'h00c8,16'h0001,-16'h0016,-16'h0021,16'h0008,16'h00da,16'h0078,16'h004d,16'h0016,-16'h0057,-16'h0041,16'h0015,-16'h0027,16'h000d,16'h0091,16'h0000,16'h0003,16'h005c,16'h003a,-16'h0009,16'h0017,16'h0007,-16'h0019,16'h0033,-16'h001d,16'h0032,16'h0010,16'h000b,16'h0058,16'h0000,16'h0057,-16'h001b,-16'h0061,-16'h0029,-16'h0013,16'h0023,-16'h0025,16'h0023,16'h003e,16'h0028,16'h0059,16'h0076,-16'h0064,16'h0016,16'h0015,-16'h0009,16'h000f,16'h002a,16'h0050,16'h0091,-16'h005a,16'h0031,16'h0000,16'h0025,16'h0000,16'h002d,-16'h003d,16'h0028,-16'h0030,-16'h000b,-16'h001f,-16'h0003,16'h001d,16'h000a,-16'h00f1,-16'h0011,-16'h0019,-16'h0029,-16'h001f,16'h00d9,16'h0061,16'h003c,16'h0003,-16'h0053,-16'h000e,-16'h0023,-16'h004b,16'h000c,16'h008f,-16'h002a,-16'h0019,16'h0061,16'h003b,-16'h0014,16'h0005,16'h0031,-16'h0010,16'h000d,-16'h0048,16'h002b,-16'h000b,-16'h001b,16'h0055,16'h0032,16'h007a,-16'h0006,-16'h0049,-16'h0032,16'h0007,16'h0015,-16'h002e,16'h0039,16'h002d,16'h0029,16'h0073,16'h0079,-16'h00a2,16'h0019,16'h0016,-16'h001c,-16'h0001,16'h0014,16'h0052,16'h0065,-16'h0099,16'h0012,-16'h0024,16'h0032,-16'h001e,16'h002f,-16'h004b,16'h0010,-16'h0016,-16'h0015,-16'h007d,-16'h0012,16'h005b,16'h002b,-16'h00db,-16'h0003,-16'h0042,-16'h0009,-16'h0021,16'h008c,16'h0035,16'h001a,-16'h002d,-16'h000d,16'h0025,-16'h006f,-16'h0034,-16'h0014,16'h0060,-16'h003e,16'h0011,16'h004b,16'h004c,-16'h001b,-16'h0013,16'h0022,16'h001a,16'h0010,-16'h002d,16'h0029,16'h001f,-16'h0034,16'h0047,16'h008a,16'h0063,-16'h000c,-16'h0040,-16'h003a,16'h0014,16'h001a,-16'h002f,16'h003f,16'h003c,16'h002c,16'h004c,16'h0066,-16'h00e1,16'h0051,16'h002b,16'h000f,16'h001d,16'h0012,16'h005c,16'h0034,-16'h009c,-16'h0008,-16'h0038,-16'h0012,-16'h0024,16'h0007,-16'h0026,16'h0011,-16'h001e,16'h001e,-16'h00b1,16'h0006,16'h007e,16'h003b,-16'h006b,16'h0046,-16'h003e,16'h0000,-16'h0016,16'h0076,16'h001b,16'h002e,-16'h006d,16'h0057,16'h000f,-16'h007a,-16'h0038,-16'h0003,16'h0079,-16'h001f,16'h000d,16'h0023,16'h0062,16'h001f,-16'h0012,16'h003b,16'h001c,16'h0029,-16'h0044,16'h002d,-16'h0008,-16'h0022,16'h004e,16'h007a,16'h002c,-16'h004d,-16'h004d,-16'h0042,16'h0018,16'h000d,-16'h006d,16'h002f,16'h001b,16'h001a,16'h0060,16'h0074,-16'h00ba,16'h006c,16'h0026,16'h0017,16'h0018,-16'h0006,16'h005e,16'h0014,-16'h006a,16'h0002,16'h0029,-16'h0046,-16'h000b,-16'h000d,-16'h0019,16'h0018,-16'h0030,16'h004b,-16'h0081,16'h001b,16'h00a0,16'h0058,-16'h0041,16'h0021,-16'h0047,16'h0002,-16'h0010,16'h008e,16'h0014,16'h0028,-16'h0052,16'h006e,-16'h0021,-16'h0087,-16'h0037,-16'h0011,16'h003a,-16'h0050,16'h0003,16'h0018,16'h0066,-16'h0002,-16'h0029,16'h0035,16'h0015,16'h0012,-16'h0024,16'h001a,-16'h0006,16'h0008,16'h003a,16'h0081,-16'h0005,-16'h0069,-16'h0067,-16'h0048,16'h0010,16'h002d,-16'h0051,16'h0044,16'h0021,-16'h000b,16'h0043,16'h0070,-16'h00b8,16'h004c,16'h0033,16'h002b,16'h003c,16'h0000,16'h005d,16'h001a,-16'h0050,16'h0025,16'h0022,16'h0001,16'h0012,16'h0004,-16'h0004,-16'h0012,-16'h0027,16'h0037,-16'h0024,16'h0042,16'h00be,16'h007a,-16'h0051,16'h0044,-16'h004d,-16'h0025,16'h001a,16'h008b,16'h002f,16'h0044,-16'h0033,16'h003f,-16'h0065,-16'h0062,-16'h0005,-16'h001f,16'h0007,-16'h002f,-16'h0035,-16'h0006,16'h0079,-16'h0002,-16'h0021,16'h004a,16'h002a,16'h0020,-16'h0024,16'h004b,-16'h0009,-16'h0005,16'h002a,16'h0058,-16'h004e,-16'h0048,-16'h007a,-16'h0045,-16'h000d,16'h001f,-16'h0062,16'h0025,16'h002d,16'h000b,16'h0053,16'h0053,-16'h00d5,16'h0040,16'h004d,16'h0036,16'h0025,16'h0019,16'h0062,16'h002e,-16'h001a,16'h0036,16'h0012,16'h0005,16'h0009,16'h0009,16'h0019,-16'h0018,-16'h0009,16'h002b,16'h0000,16'h003f,16'h00a1,16'h006b,-16'h005e,16'h0047,-16'h002a,-16'h006c,16'h0021,16'h007d,16'h0060,16'h002c,16'h001b,-16'h0027,-16'h005c,-16'h0018,16'h003b,-16'h0021,-16'h0020,16'h0027,-16'h005c,-16'h0002,16'h006e,-16'h000a,-16'h0011,16'h0022,16'h002c,16'h002e,-16'h0020,16'h0050,-16'h0011,16'h0036,-16'h000e,16'h0061,-16'h006e,-16'h001a,-16'h006b,16'h000e,16'h0001,16'h0050,-16'h003b,-16'h0002,-16'h0007,16'h000a,16'h005f,16'h0052,-16'h00e7,16'h003a,16'h004d,16'h0028,16'h0032,16'h0002,16'h005e,16'h0051,16'h0023,16'h0042,-16'h0009,16'h004f,16'h0000,16'h0012,16'h002b,-16'h003a,-16'h0008,-16'h0019,16'h0019,16'h003b,16'h0072,16'h0019,-16'h0070,16'h0025,-16'h002b,-16'h0066,-16'h0002,16'h006b,16'h005c,16'h0031,16'h001a,-16'h0050,16'h000e,-16'h0005,16'h0037,16'h0009,-16'h0016,16'h0037,-16'h0081,-16'h001a,16'h0060,16'h000f,-16'h0013,16'h0026,-16'h0004,16'h0022,-16'h0030,16'h0020,-16'h0016,16'h0031,-16'h001c,16'h003f,-16'h0060,16'h0003,-16'h0092,16'h0017,16'h0005,16'h004d,-16'h0021,-16'h002b,16'h002e,-16'h0016,16'h006d,16'h002a,-16'h00b7,16'h004e,16'h002f,16'h0034,16'h003e,16'h0029,16'h003e,16'h005a,16'h003d,16'h0037,-16'h003b,16'h0037,16'h000e,-16'h0027,16'h0030,-16'h0028,16'h0007,-16'h0013,16'h0048,16'h003b,16'h0098,-16'h0085,-16'h0052,-16'h0017,16'h0001,-16'h0008,16'h001d,16'h0026,16'h0048,16'h0031,16'h003e,-16'h0032,16'h0051,16'h0016,-16'h0047,16'h001e,-16'h000d,16'h0038,-16'h004f,-16'h0012,16'h006c,16'h0021,-16'h0001,16'h001d,-16'h0007,16'h0003,-16'h001d,16'h0030,16'h0005,16'h0039,-16'h0055,16'h0013,-16'h0001,-16'h0008,-16'h0080,16'h0029,16'h0037,16'h0060,-16'h003e,16'h0000,16'h002a,-16'h0029,16'h0075,16'h0028,-16'h0091,16'h004c,16'h0039,16'h002b,16'h000c,16'h0000,16'h0045,16'h002a,16'h0045,16'h0043,-16'h003a,16'h0036,16'h0012,-16'h0049,16'h0033,-16'h001f,16'h000e,-16'h0011,16'h0054,16'h0005,16'h0096,-16'h0082,-16'h004e,-16'h0001,-16'h000d,16'h0050,16'h003a,-16'h0039,16'h0007,16'h0036,16'h001b,16'h000a,16'h0027,16'h0024,-16'h0090,-16'h0015,16'h0011,16'h0042,-16'h003e,-16'h0016,16'h004e,16'h0036,16'h0003,16'h001d,16'h0004,16'h0008,-16'h0021,16'h0050,-16'h0010,16'h0034,-16'h0035,-16'h000c,16'h0027,16'h0027,-16'h001f,16'h0029,16'h0039,16'h0037,-16'h0023,-16'h0005,16'h0005,-16'h000e,16'h000c,16'h0025,-16'h0087,16'h0049,16'h001d,-16'h0006,16'h000d,16'h000d,16'h0037,16'h002a,16'h004d,16'h0066,-16'h002b,16'h001e,16'h001b,-16'h0020,16'h0055,-16'h000c,16'h0012,16'h0001,16'h0030,-16'h0014,16'h0074,-16'h0083,-16'h0065,16'h0004,-16'h001f,16'h0074,16'h0028,-16'h005d,-16'h0081,16'h0046,16'h0015,16'h004e,16'h0005,-16'h0007,-16'h0080,-16'h001d,-16'h0012,16'h002b,-16'h0014,-16'h0008,16'h0034,16'h003a,-16'h0005,16'h0043,16'h0008,-16'h0006,-16'h0033,16'h0072,-16'h0013,16'h0019,-16'h002c,16'h000d,16'h0076,16'h0018,-16'h0010,16'h0046,16'h0013,16'h000a,-16'h0025,-16'h0017,16'h002d,-16'h000a,-16'h000c,16'h001f,-16'h0075,16'h0050,16'h001a,-16'h0014,16'h001f,16'h000f,16'h004d,16'h0000,16'h0038,16'h0031,-16'h0007,16'h000a,-16'h000f,16'h0020,16'h005d,16'h0010,16'h000b,16'h0032,16'h0015,-16'h0012,16'h0095,-16'h0051,-16'h0083,-16'h0010,-16'h0042,16'h0070,16'h000c,-16'h005c,-16'h0087,16'h0037,16'h0004,16'h0027,-16'h0013,-16'h0004,-16'h003c,-16'h0002,-16'h001c,16'h0007,16'h0020,-16'h0003,16'h0023,16'h002e,16'h0022,16'h0036,16'h001f,-16'h0024,-16'h0004,16'h006b,-16'h001b,-16'h000a,-16'h0032,-16'h0011,16'h0082,-16'h0008,-16'h0014,16'h0043,16'h000a,16'h0011,-16'h002d,-16'h0018,16'h0012,-16'h001a,16'h000b,16'h0012,-16'h0069,16'h0029,16'h0015,-16'h0033,16'h0034,-16'h0010,16'h0040,16'h001b,16'h003f,16'h0041,-16'h0004,-16'h000c,-16'h0006,16'h0001,16'h004f,16'h0006,16'h001b,16'h0026,-16'h0018,-16'h0016,16'h006e,-16'h0038,-16'h0076,-16'h000b,-16'h002a,16'h0037,-16'h001e,-16'h0061,-16'h00a6,16'h0036,16'h0020,16'h0021,16'h0029,-16'h001c,16'h0018,-16'h0016,16'h0029,16'h0032,16'h0000,16'h000e,16'h0008,16'h001b,16'h000d,16'h004d,16'h0002,16'h0006,-16'h000e,16'h0065,-16'h0007,16'h000f,-16'h005b,-16'h0001,16'h006a,-16'h000a,16'h0005,16'h0027,16'h001f,16'h0007,16'h0004,-16'h0024,16'h0024,-16'h0013,16'h002b,16'h0019,-16'h0052,16'h002b,16'h0020,-16'h005a,16'h0010,-16'h0050,16'h0062,16'h001e,16'h004d,16'h0064,-16'h0007,-16'h0014,16'h0024,-16'h000c,16'h0061,16'h0013,16'h0032,16'h002f,-16'h0019,16'h0007,16'h006a,16'h001e,-16'h006f,16'h0045,-16'h001f,16'h001d,-16'h0009,-16'h0032,-16'h0069,16'h0037,16'h0044,16'h0007,16'h0055,-16'h0027,16'h0055,-16'h0024,16'h002d,16'h002d,-16'h0016,-16'h000c,16'h000b,16'h004d,16'h0003,16'h0051,16'h0017,16'h0023,-16'h0009,16'h005c,16'h000f,16'h001e,-16'h0035,-16'h002c,-16'h004d,-16'h001f,16'h001e,16'h0031,16'h0023,16'h000e,-16'h0027,-16'h0042,16'h0017,16'h0016,16'h0062,16'h0027,-16'h0070,16'h001e,16'h0008,-16'h0049,-16'h0011,-16'h0097,16'h0023,16'h0038,16'h002e,16'h0066,-16'h001d,-16'h001d,16'h0000,-16'h002a,16'h004e,-16'h0009,16'h0015,16'h003a,-16'h0015,-16'h000d,16'h0050,16'h002c,-16'h0043,16'h003b,-16'h0001,-16'h0016,-16'h002e,-16'h000e,-16'h0046,16'h004b,16'h0030,-16'h0048,16'h0029,-16'h0021,16'h0032,-16'h001e,16'h0020,16'h0025,-16'h0029,16'h000f,-16'h000f,16'h005b,-16'h0003,16'h003b,16'h0017,16'h0038,-16'h0028,16'h006a,-16'h0007,16'h001d,-16'h0014,-16'h0053,-16'h008b,-16'h002b,16'h0046,16'h001a,16'h0046,16'h000b,-16'h001b,-16'h0020,16'h001f,16'h0033,16'h0085,16'h000c,-16'h0085,16'h0000,16'h001b,-16'h0046,-16'h0024,-16'h00d8,16'h002a,16'h0023,16'h0008,16'h004a,-16'h0014,-16'h000a,-16'h0005,-16'h0019,16'h0062,16'h000d,16'h0014,16'h0027,-16'h001f,16'h001b,16'h004f,16'h0011,16'h0002,16'h0051,16'h0016,-16'h0034,-16'h0037,-16'h0008,-16'h001c,16'h0057,16'h002f,-16'h004c,-16'h0003,-16'h0039,16'h001f,-16'h0017,16'h0030,16'h0021,-16'h0017,16'h0024,-16'h0012,16'h0037,-16'h0006,16'h0019,16'h0043,16'h0037,-16'h002b,16'h0064,-16'h0015,16'h0053,16'h0004,-16'h003b,-16'h00ae,-16'h0014,16'h0044,-16'h000f,16'h002d,16'h0032,-16'h0029,-16'h0012,16'h0031,16'h0005,16'h0082,16'h0028,-16'h0063,-16'h0003,16'h0022,-16'h0038,16'h0010,-16'h0132,16'h001a,16'h0038,16'h0014,16'h005d,-16'h0031,-16'h0010,16'h0003,16'h000d,16'h0051,16'h000c,16'h0027,16'h001c,-16'h0008,16'h003a,16'h003e,16'h0040,-16'h003e,16'h0070,16'h0010,16'h0012,16'h0006,-16'h004c,16'h001f,16'h0045,16'h0019,-16'h0044,-16'h000d,-16'h0032,16'h0001,16'h000a,16'h0067,16'h004c,16'h004e,16'h001f,16'h000f,16'h000d,-16'h0044,16'h0039,16'h0016,16'h0053,-16'h0001,16'h006c,-16'h0035,16'h0023,16'h0002,-16'h0054,-16'h0060,-16'h0011,16'h0035,-16'h0015,16'h0065,16'h0049,-16'h002d,-16'h001b,16'h005e,16'h0018,16'h0083,16'h0022,-16'h006a,16'h0006,16'h003d,-16'h0046,16'h0018,-16'h0181,16'h000b,16'h0011,16'h0016,16'h0052,-16'h000f,16'h0002,-16'h001b,-16'h0003,16'h004f,-16'h0011,16'h0006,16'h0029,-16'h0002,16'h0033,16'h0048,16'h0041,-16'h0013,16'h0065,16'h002c,16'h0010,16'h0033,-16'h003a,16'h0012,16'h0057,16'h0006,-16'h0008,-16'h0052,-16'h0009,-16'h0015,-16'h001d,16'h0022,16'h001d,16'h0060,16'h0037,16'h0038,-16'h0007,-16'h002e,16'h0067,16'h001c,16'h0043,-16'h001b,16'h0049,-16'h001e,16'h0052,-16'h0005,-16'h0069,16'h0018,-16'h002b,16'h002c,-16'h0024,16'h0057,16'h003f,-16'h0063,-16'h0023,16'h0036,16'h0004,16'h0052,16'h0036,-16'h0044,16'h0039,16'h003a,-16'h0032,16'h005c,-16'h01fe,16'h0025,16'h000e,16'h001c,16'h0052,-16'h0022,16'h000c,-16'h000a,16'h0009,16'h003e,-16'h0003,-16'h0017,-16'h0009,-16'h000a,16'h000a,16'h0041,16'h0029,-16'h001b,16'h0025,16'h0032,16'h001e,16'h0058,-16'h003c,16'h000d,16'h005e,-16'h0010,16'h0019,-16'h0026,16'h0016,-16'h003e,-16'h0026,16'h0024,16'h0021,16'h0045,16'h002d,16'h0031,16'h0018,-16'h005e,16'h005b,16'h0010,16'h002f,-16'h001d,16'h0041,-16'h0029,16'h003a,-16'h0016,-16'h0055,16'h005b,-16'h0015,16'h0040,-16'h0009,16'h0038,16'h004b,-16'h0071,16'h0019,16'h002d,16'h0026,16'h003f,16'h0020,-16'h0048,16'h0033,16'h002d,-16'h002d,16'h003a,-16'h0200,16'h000f,-16'h0010,-16'h0012,16'h005b,-16'h001e,16'h003b,16'h002f,16'h0029,16'h0036,16'h0017,-16'h0004,16'h0059,16'h0011,-16'h0012,16'h003b,16'h0022,-16'h0005,-16'h00bc,16'h0048,-16'h0005,16'h005b,-16'h0020,16'h0021,16'h0066,-16'h000a,16'h0056,-16'h003f,16'h0001,-16'h003c,-16'h003c,16'h0006,16'h0011,16'h0017,16'h0048,16'h0045,16'h001c,-16'h00b4,16'h0049,-16'h000a,16'h0026,-16'h0031,16'h003f,16'h000e,16'h0007,-16'h0018,-16'h003d,16'h0039,-16'h0001,16'h0032,-16'h0011,16'h0019,16'h0025,-16'h006f,-16'h0002,16'h000d,-16'h0005,16'h0001,-16'h001c,-16'h0044,16'h005f,16'h0009,-16'h0011,16'h0026,-16'h01cd,16'h001b,16'h0018,16'h001b,16'h0045,16'h0009,16'h0032,16'h000f,16'h001c,16'h0025,16'h0027,16'h0015,16'h0012,-16'h0001,-16'h004c,16'h0048,16'h0010,-16'h0017,-16'h023d,16'h004c,16'h0002,16'h0075,-16'h0051,16'h001a,16'h0061,16'h0008,16'h006a,-16'h0022,16'h001f,-16'h002a,-16'h003a,16'h000e,16'h0001,16'h0000,16'h0037,16'h0026,16'h003c,-16'h00f2,16'h004e,-16'h0032,16'h001b,-16'h0030,16'h0054,16'h000a,-16'h0026,-16'h0030,-16'h002b,16'h0014,16'h0012,16'h0018,-16'h002f,-16'h0080,16'h0008,-16'h0059,-16'h000e,16'h0016,-16'h001c,16'h0032,-16'h0015,-16'h0030,16'h006c,16'h0011,-16'h000f,16'h002a,-16'h0154,16'h000a,16'h0013,16'h001d,16'h001c,16'h0028,16'h0008,16'h0031,16'h0008,16'h0046,16'h000a,16'h0034,-16'h007a,-16'h0028,-16'h0092,16'h005f,-16'h0020,-16'h0045,-16'h02ac,16'h005e,16'h0028,16'h008b,-16'h005f,-16'h0010,16'h003e,16'h0059,16'h0079,-16'h003c,16'h0005,-16'h0012,-16'h0058,16'h0018,16'h0021,16'h0013,16'h0038,-16'h000c,16'h0009,-16'h00c4,16'h002a,-16'h002d,16'h0035,-16'h0037,16'h0066,16'h0016,16'h0008,-16'h002d,16'h0002,-16'h0022,16'h0027,16'h0069,-16'h000e,-16'h01e3,16'h0021,-16'h0074,-16'h0018,16'h0027,-16'h0051,16'h0055,16'h0009,-16'h001e,16'h0057,-16'h0016,16'h0006,16'h0021,-16'h010f,16'h0039,16'h0031,16'h0020,16'h0014,16'h002f,-16'h0013,16'h0007,-16'h000b,16'h004e,16'h0036,16'h0007,-16'h00b7,-16'h001a,-16'h00d3,16'h002e,-16'h003a,-16'h003c,-16'h0156,16'h005e,16'h0037,16'h003e,-16'h007c,-16'h0034,16'h0049,16'h0027,16'h004a,16'h0000,16'h0002,16'h0037,-16'h0036,16'h0012,16'h0023,16'h0021,16'h004b,16'h000e,16'h0005,-16'h00c6,16'h0032,-16'h003f,16'h0018,16'h000a,16'h0055,16'h0003,16'h0022,16'h000f,16'h000e,-16'h001e,16'h0008,16'h003f,-16'h002f,-16'h022e,16'h0019,-16'h004f,16'h0002,16'h0004,-16'h0072,16'h005f,16'h000c,-16'h0018,16'h0057,-16'h000f,-16'h0016,16'h001b,-16'h00c3,16'h0017,16'h0067,16'h000f,16'h000f,16'h0047,-16'h0023,-16'h0015,-16'h0003,16'h002f,-16'h0003,-16'h0002,-16'h008a,-16'h0025,-16'h0103,16'h004d,-16'h0046,-16'h0028,-16'h00c0,16'h0063,16'h0007,-16'h00d5,-16'h005b,-16'h0065,16'h0052,-16'h0017,16'h006a,16'h0029,-16'h0009,16'h0047,-16'h0037,16'h003f,16'h0015,16'h0006,16'h006e,-16'h0003,16'h0017,-16'h00d4,16'h000f,-16'h0046,-16'h0017,16'h003e,16'h0045,16'h001a,16'h0026,16'h0045,16'h0011,16'h0014,16'h0004,16'h003c,16'h0000,-16'h012d,16'h003e,-16'h004c,-16'h002b,16'h0017,-16'h005c,16'h005a,16'h0011,-16'h0006,16'h003a,-16'h001a,-16'h0041,-16'h003b,-16'h00af,16'h0035,16'h0099,16'h002e,-16'h0011,16'h0028,-16'h0014,-16'h0027,16'h0014,16'h004a,-16'h0018,16'h0001,-16'h007e,-16'h0004,-16'h00d5,16'h003a,-16'h0016,-16'h003c,-16'h005b,16'h006e,16'h0018,-16'h01a0,-16'h003b,-16'h00b0,16'h0014,-16'h0004,16'h0075,16'h0011,16'h000b,16'h002e,-16'h0046,16'h0029,-16'h0001,-16'h0001,16'h0087,-16'h0006,-16'h0002,-16'h00bd,16'h0003,-16'h004a,-16'h0007,16'h0094,16'h003e,16'h0054,16'h0038,16'h007e,-16'h0018,-16'h000c,-16'h0028,16'h0032,16'h0004,-16'h007c,16'h0045,-16'h0071,-16'h0039,16'h0019,-16'h0024,16'h0064,16'h0028,-16'h0004,-16'h001e,-16'h001e,-16'h002f,-16'h0048,-16'h008d,16'h0017,16'h00a1,16'h0014,-16'h005d,16'h0053,-16'h0003,-16'h004f,16'h001d,16'h0069,-16'h001a,16'h0020,-16'h0051,-16'h0030,-16'h0087,16'h002d,-16'h0015,-16'h0036,-16'h0009,16'h0088,16'h0021,-16'h0194,-16'h000c,-16'h00a3,16'h0019,-16'h0041,16'h003c,16'h0022,16'h0011,16'h001d,-16'h000c,16'h002d,-16'h0001,16'h0001,16'h0045,16'h0034,16'h0027,-16'h0090,-16'h0033,-16'h000a,-16'h0003,16'h0099,16'h0041,16'h005d,16'h0033,16'h00a0,16'h000e,-16'h0006,-16'h000d,16'h003a,-16'h0004,-16'h0029,-16'h0017,-16'h0034,-16'h0011,16'h0003,-16'h000b,16'h0061,16'h0000,-16'h0003,-16'h0078,-16'h0034,-16'h0003,-16'h004e,-16'h00a0,-16'h0022,16'h0089,16'h0021,-16'h000f,16'h0022,16'h0034,-16'h006e,16'h004b,16'h0070,-16'h001b,16'h002b,-16'h0039,-16'h0022,-16'h004e,16'h0031,-16'h001d,-16'h0032,16'h0028,16'h007d,16'h0037,-16'h00ef,-16'h0012,-16'h0093,16'h0028,-16'h004c,-16'h0009,16'h0003,16'h0032,16'h0012,16'h0005,16'h0023,16'h0003,16'h005d,16'h0041,16'h005e,16'h0011,-16'h0093,-16'h000d,-16'h0025,-16'h001c,16'h004f,16'h005a,16'h0019,16'h0000,16'h0081,16'h0005,-16'h0014,-16'h0024,16'h001d,16'h0015,16'h0004,-16'h004e,-16'h0041,16'h0035,16'h004c,16'h0026,16'h002f,16'h0035,-16'h0050,16'h0022,16'h0043,16'h0011,16'h003f,16'h0060,-16'h001d,16'h009b,-16'h0032,16'h0095,-16'h0009,-16'h0004,16'h0026,16'h0008,16'h000a,16'h0009,-16'h0059,-16'h004d,16'h000e,16'h007e,-16'h0030,-16'h002b,-16'h0087,16'h0016,-16'h0015,16'h0021,-16'h0008,16'h00c8,16'h0066,16'h004c,16'h0028,-16'h0056,-16'h001b,16'h0060,-16'h0015,-16'h0018,16'h0078,16'h0008,16'h0014,16'h0020,16'h0009,16'h0015,-16'h0006,16'h000b,16'h003b,16'h0025,-16'h0018,16'h0082,-16'h0011,16'h0014,16'h002e,-16'h0024,16'h0016,-16'h002b,-16'h0046,-16'h003f,-16'h0022,16'h0083,-16'h0010,16'h004e,16'h0039,16'h0037,16'h0037,16'h0024,-16'h0063,16'h0039,16'h0031,16'h0019,16'h0045,16'h004c,16'h0001,16'h009c,-16'h0054,16'h007d,-16'h0004,16'h0006,16'h0026,16'h0028,-16'h000f,16'h000c,-16'h005b,-16'h0025,16'h000d,16'h0040,16'h000d,-16'h0005,-16'h00c3,16'h000b,16'h000a,16'h002c,-16'h0030,16'h00e1,16'h0077,16'h0019,16'h0008,-16'h0044,-16'h0022,16'h003d,-16'h0017,-16'h001b,16'h0086,-16'h0008,16'h000a,16'h001e,16'h0023,-16'h000c,16'h000c,-16'h0007,16'h0005,16'h0020,-16'h0026,16'h0059,16'h0000,16'h001e,16'h0049,16'h0025,16'h005b,-16'h000f,-16'h0058,-16'h005c,-16'h0036,16'h004a,16'h0007,16'h0043,16'h0044,16'h0032,16'h0034,16'h0035,-16'h007e,16'h0048,16'h002f,-16'h0009,16'h001a,16'h002a,16'h0059,16'h00a3,-16'h0092,16'h0061,-16'h0002,16'h0021,-16'h0002,16'h003a,-16'h0021,-16'h0020,-16'h004f,-16'h002f,16'h000a,16'h000e,-16'h0014,16'h0000,-16'h00f0,-16'h001b,-16'h0027,16'h0000,-16'h000f,16'h00c4,16'h0090,16'h0042,-16'h0005,-16'h0058,-16'h0013,-16'h0021,-16'h0040,-16'h000b,16'h009a,-16'h0020,-16'h0035,16'h0005,16'h0040,-16'h0006,16'h0017,16'h002e,16'h000a,16'h001d,-16'h003c,16'h0033,16'h0000,16'h0004,16'h0087,16'h0057,16'h0077,16'h0007,-16'h0045,-16'h0062,-16'h0001,16'h0010,-16'h000f,16'h003e,16'h0034,16'h0028,16'h0053,16'h002f,-16'h0075,16'h0058,16'h0047,-16'h0002,16'h0003,16'h0019,16'h007f,16'h0068,-16'h0058,-16'h0001,16'h0007,16'h0018,-16'h0021,16'h0008,-16'h0043,-16'h0036,-16'h002c,-16'h0011,-16'h0045,16'h0000,16'h0033,16'h002d,-16'h00ce,16'h0000,-16'h003a,-16'h0001,-16'h0034,16'h009d,16'h0057,16'h000c,-16'h002b,-16'h0008,16'h0000,-16'h0040,-16'h0028,-16'h0018,16'h0082,-16'h0037,-16'h0009,16'h0024,16'h0031,-16'h0009,16'h0004,16'h001a,16'h001a,16'h002a,-16'h003e,16'h0017,16'h0005,-16'h0020,16'h0064,16'h0077,16'h0047,-16'h0007,-16'h0027,-16'h0053,16'h0001,16'h0001,-16'h0032,16'h0073,16'h000d,16'h004b,16'h005b,16'h004b,-16'h0080,16'h0083,16'h0025,16'h0006,16'h0007,16'h0007,16'h007d,16'h0047,-16'h0043,-16'h0039,16'h0008,16'h0006,-16'h002a,16'h0017,-16'h0069,-16'h0006,-16'h0013,16'h0008,-16'h0081,-16'h0003,16'h006a,16'h004c,-16'h006b,16'h002b,-16'h0051,16'h0028,-16'h0002,16'h005e,16'h0042,16'h0004,-16'h002f,16'h0010,16'h0003,-16'h0047,-16'h002d,-16'h0033,16'h008d,-16'h0051,16'h000a,16'h0019,16'h0021,-16'h0009,16'h000a,16'h001b,16'h001b,16'h002a,-16'h006c,16'h0017,-16'h001d,-16'h000c,16'h006e,16'h0062,16'h0015,-16'h0035,-16'h0056,-16'h0052,16'h0017,16'h003b,-16'h0047,16'h0062,-16'h0008,16'h002e,16'h0060,16'h005d,-16'h0064,16'h008c,16'h0048,16'h002e,-16'h0009,-16'h0001,16'h0090,16'h0034,-16'h004f,-16'h0056,16'h0015,-16'h0021,-16'h002c,16'h0006,-16'h007b,-16'h001b,-16'h0019,16'h0027,-16'h0072,-16'h0017,16'h0074,16'h0084,-16'h0004,16'h000d,-16'h004d,-16'h0015,16'h0010,16'h0073,16'h0039,16'h0030,-16'h0037,16'h0049,-16'h0024,-16'h0083,-16'h0038,-16'h0028,16'h0089,-16'h003c,-16'h0011,16'h000d,16'h004a,-16'h0008,16'h0000,16'h0036,16'h0002,-16'h0001,-16'h0023,16'h001e,-16'h0015,-16'h001f,16'h0044,16'h0085,-16'h000a,-16'h0044,-16'h0065,-16'h003d,-16'h0006,16'h002a,-16'h0054,16'h005e,16'h0007,16'h0012,16'h0055,16'h0052,-16'h0061,16'h0091,16'h003e,16'h0031,16'h0018,-16'h0006,16'h0084,16'h003a,-16'h0041,-16'h003a,16'h001f,-16'h002d,16'h0006,16'h001d,-16'h005f,-16'h0021,-16'h0016,16'h0042,-16'h003a,16'h0023,16'h0082,16'h0059,-16'h0046,16'h0022,-16'h0050,-16'h0035,16'h0035,16'h006f,16'h002f,16'h0026,-16'h000b,16'h002e,-16'h0066,-16'h0047,16'h0035,-16'h0028,16'h0052,-16'h001e,-16'h0025,16'h0001,16'h0040,16'h0004,-16'h0009,16'h002c,-16'h0009,16'h0019,-16'h0011,16'h0023,-16'h002f,-16'h0027,16'h001f,16'h0042,-16'h0051,-16'h0040,-16'h0051,-16'h0027,16'h0000,16'h0049,-16'h0045,16'h0043,-16'h0018,16'h0013,16'h005c,16'h001a,-16'h006a,16'h0092,16'h004c,16'h004b,16'h001c,16'h000d,16'h0097,16'h002c,16'h0004,-16'h0031,16'h0018,16'h0004,16'h0019,16'h0051,-16'h001f,-16'h0045,-16'h000e,16'h0048,16'h0002,16'h0027,16'h008f,16'h004d,-16'h0055,-16'h0008,-16'h0041,-16'h0048,16'h0027,16'h0052,16'h002a,16'h0033,16'h002e,-16'h0034,-16'h004b,-16'h0023,16'h003f,-16'h0017,16'h0054,16'h000c,-16'h0050,-16'h0009,16'h003e,16'h0005,-16'h0012,16'h0029,16'h0017,16'h0031,16'h000b,16'h001d,-16'h002a,16'h0006,16'h0008,16'h002d,-16'h0053,-16'h0008,-16'h0076,-16'h000b,-16'h0003,16'h004d,-16'h0057,16'h0019,-16'h0021,16'h0003,16'h0053,-16'h000a,-16'h0067,16'h006d,16'h0056,16'h001d,16'h001c,16'h0015,16'h008b,16'h003b,16'h003d,-16'h003e,-16'h0005,16'h0020,16'h0019,16'h003c,16'h000f,-16'h003c,16'h000c,16'h000c,-16'h0001,16'h0020,16'h0072,16'h000d,-16'h0065,16'h0011,-16'h0038,-16'h0070,16'h0005,16'h0076,16'h0032,16'h0023,16'h0054,-16'h0072,16'h0004,16'h001b,16'h002b,16'h0007,16'h002c,16'h0006,-16'h004f,-16'h001c,16'h003b,16'h002a,-16'h001f,16'h001a,-16'h0012,16'h001f,16'h000f,-16'h001d,-16'h0023,16'h001e,-16'h0024,16'h0016,-16'h0031,16'h0010,-16'h009d,16'h000f,16'h0017,16'h0043,-16'h0029,16'h000f,-16'h0004,-16'h001f,16'h006c,-16'h003f,-16'h0081,16'h0080,16'h0026,16'h0004,16'h0023,-16'h0016,16'h0079,16'h0018,16'h0053,-16'h0011,-16'h0033,16'h002c,16'h0029,-16'h0003,16'h002c,-16'h0043,16'h0012,-16'h0027,16'h0005,16'h0007,16'h0092,-16'h0059,-16'h0039,16'h0000,-16'h0045,-16'h0030,16'h0036,16'h0061,16'h0033,16'h002d,16'h0011,-16'h002d,16'h0018,16'h0039,-16'h0051,16'h0000,16'h0028,-16'h000b,-16'h0051,-16'h0050,16'h0037,-16'h0010,-16'h000d,16'h000b,16'h000c,16'h0025,-16'h0008,-16'h0002,-16'h0026,16'h003e,-16'h0044,-16'h0006,-16'h0010,16'h0019,-16'h007a,16'h0024,16'h0033,16'h004e,-16'h0038,16'h0011,-16'h001d,-16'h0014,16'h0067,-16'h002c,-16'h004d,16'h00ac,16'h0030,16'h000b,16'h001f,-16'h0025,16'h0095,16'h0028,16'h003f,-16'h0005,-16'h0041,16'h0037,16'h000f,16'h0012,16'h003d,16'h0000,-16'h000a,-16'h000e,16'h000b,16'h0004,16'h0087,-16'h005d,-16'h0023,-16'h000c,-16'h004c,16'h002a,16'h004c,16'h004a,-16'h0032,16'h002e,16'h0035,16'h0010,16'h0020,16'h001d,-16'h00ae,-16'h0009,16'h0030,16'h0018,-16'h0047,-16'h0032,16'h001c,16'h0025,16'h0004,16'h0045,16'h0004,16'h0022,-16'h001e,16'h000c,-16'h000f,16'h0051,-16'h0038,-16'h0014,16'h0030,16'h0020,-16'h0078,16'h0019,16'h004b,16'h002e,-16'h0042,16'h0005,-16'h0046,-16'h001a,16'h0047,16'h000d,-16'h0081,16'h00a8,16'h0010,-16'h0026,16'h0018,-16'h0063,16'h008e,16'h0022,16'h0053,-16'h000c,-16'h002d,16'h0025,16'h0016,16'h0026,16'h0053,-16'h000b,-16'h0002,16'h0007,16'h0026,16'h000d,16'h0096,-16'h0041,-16'h0016,-16'h000d,-16'h005a,16'h0066,16'h0018,16'h002e,-16'h0079,16'h0049,16'h0016,16'h0034,-16'h002f,16'h0000,-16'h008b,-16'h0035,16'h0038,-16'h0014,-16'h0009,-16'h002d,-16'h0009,16'h0026,-16'h002b,16'h0041,16'h0002,16'h0021,-16'h0033,16'h0035,-16'h002a,16'h0013,-16'h0004,16'h0005,16'h0044,16'h0023,-16'h0084,16'h0012,16'h004a,16'h002a,-16'h0042,-16'h0013,-16'h002d,16'h0018,16'h0013,16'h000c,-16'h006d,16'h00b9,16'h0000,-16'h0039,16'h002f,-16'h009a,16'h0072,16'h000b,16'h004b,-16'h002d,-16'h000a,16'h001f,16'h000b,16'h0044,16'h005a,-16'h0002,-16'h000b,16'h0013,-16'h0007,16'h000a,16'h0095,-16'h004f,-16'h0066,-16'h0004,-16'h0071,16'h005a,-16'h0003,16'h0029,-16'h0091,16'h0053,-16'h0002,16'h0023,-16'h001d,-16'h0017,-16'h0054,-16'h002e,16'h002c,-16'h0003,16'h000d,-16'h0041,16'h0003,16'h002e,-16'h000d,16'h0039,-16'h0005,16'h000d,-16'h002d,16'h0049,-16'h0031,16'h0023,-16'h0023,16'h0008,16'h0043,16'h0018,-16'h0048,-16'h0005,16'h0058,16'h0002,-16'h002c,-16'h0021,-16'h0027,-16'h0008,16'h0012,-16'h0026,-16'h0044,16'h00a0,16'h0000,-16'h0060,16'h0041,-16'h00bf,16'h007f,-16'h0005,16'h004c,-16'h0032,-16'h001f,16'h0000,16'h0005,16'h003b,16'h0049,-16'h000b,16'h001c,16'h0024,16'h000f,-16'h0002,16'h006d,-16'h0035,-16'h0094,16'h0001,-16'h0085,16'h0042,-16'h0011,16'h0000,-16'h0058,16'h0037,-16'h0006,16'h0000,16'h0001,-16'h004c,-16'h0021,-16'h000b,16'h0002,-16'h0022,-16'h0005,-16'h0016,-16'h0001,16'h003d,-16'h0019,16'h003f,16'h0010,16'h001b,-16'h002a,16'h0032,-16'h0048,16'h0024,-16'h001e,-16'h0017,16'h0037,-16'h000d,-16'h0015,16'h0002,16'h003a,-16'h000d,-16'h002b,-16'h002b,-16'h0005,16'h0019,16'h0016,-16'h0034,-16'h0037,16'h0065,16'h0013,-16'h0048,16'h000f,-16'h0124,16'h0082,16'h0004,16'h005b,-16'h003b,-16'h0029,-16'h001d,-16'h0010,16'h001f,16'h002d,16'h0000,16'h001d,16'h002d,16'h0006,16'h000d,16'h0053,16'h0003,-16'h0065,16'h0023,-16'h00b0,16'h003a,-16'h0004,-16'h0015,-16'h0047,16'h001f,16'h0009,-16'h0036,16'h0029,-16'h003e,16'h003e,-16'h000f,16'h0017,-16'h000f,-16'h002b,-16'h0018,-16'h0017,16'h0041,-16'h001a,16'h0037,16'h0010,16'h0036,-16'h002f,16'h005b,-16'h002d,16'h0001,-16'h0039,-16'h003e,-16'h005d,-16'h0017,16'h000d,-16'h0006,16'h002e,-16'h0011,-16'h0039,-16'h001e,16'h000f,16'h002a,16'h0043,-16'h0048,16'h0000,16'h005f,16'h0013,-16'h0035,16'h000a,-16'h0165,16'h007e,-16'h0006,16'h004f,-16'h0043,-16'h003b,-16'h0026,-16'h0015,16'h0008,16'h004f,16'h000d,16'h002a,16'h0022,16'h0006,16'h0021,16'h0069,16'h0001,-16'h0013,16'h0049,-16'h008e,16'h0014,-16'h001d,-16'h0019,-16'h001c,16'h0029,16'h0015,-16'h004c,16'h0018,-16'h0044,16'h0030,-16'h0043,16'h0022,-16'h0018,-16'h0048,-16'h0001,-16'h0007,16'h004d,-16'h0011,16'h0038,16'h001f,16'h0037,-16'h000c,16'h004d,-16'h002e,16'h0010,-16'h001a,-16'h0021,-16'h00a5,-16'h003d,16'h0013,16'h0004,16'h004e,-16'h000f,-16'h0038,-16'h002a,-16'h000e,16'h001c,16'h0061,-16'h003e,-16'h0050,16'h0045,16'h001c,-16'h002c,-16'h0022,-16'h01c6,16'h0070,-16'h0001,16'h0033,-16'h003e,-16'h0032,-16'h0028,16'h0000,16'h0005,16'h003f,16'h000f,16'h0000,16'h0016,-16'h001c,16'h0015,16'h006b,16'h000b,-16'h001c,16'h0062,-16'h0092,-16'h0044,-16'h0036,-16'h0003,-16'h0005,16'h0048,16'h003a,-16'h0073,16'h0012,-16'h0067,16'h0030,-16'h0004,16'h002a,-16'h0008,-16'h000c,16'h0027,-16'h0006,16'h0043,-16'h0052,16'h0049,16'h001c,16'h0047,-16'h001a,16'h003f,-16'h0023,16'h0018,-16'h0035,-16'h001d,-16'h00b2,-16'h0066,16'h0027,-16'h0001,16'h0053,16'h0003,-16'h002c,-16'h001f,16'h0011,16'h0001,16'h0069,-16'h0044,-16'h0038,16'h003c,16'h0037,-16'h004f,16'h0002,-16'h01ed,16'h003e,16'h000e,16'h000f,-16'h0048,-16'h002e,-16'h001b,-16'h002d,16'h0020,16'h004f,-16'h0003,16'h000b,16'h000e,-16'h0028,16'h003c,16'h0052,16'h0024,-16'h0050,16'h0059,-16'h007c,16'h0002,16'h001a,-16'h000f,-16'h0001,16'h003e,16'h0003,-16'h003c,-16'h0025,-16'h004e,-16'h0001,-16'h0009,16'h003d,16'h000e,16'h0041,16'h0039,16'h000e,16'h0016,-16'h0082,16'h004a,16'h0010,16'h004e,-16'h0029,16'h002c,-16'h0034,16'h0033,-16'h0039,-16'h0055,-16'h0040,-16'h004f,16'h0047,-16'h0012,16'h002b,16'h0024,-16'h0044,-16'h0019,-16'h0006,-16'h0008,16'h0067,16'h0018,-16'h005c,16'h002e,16'h003c,-16'h0024,16'h0019,-16'h023e,16'h001f,-16'h0013,16'h0018,-16'h0021,-16'h0015,16'h001d,-16'h000b,16'h0009,16'h0057,16'h0015,16'h0000,16'h0019,-16'h0012,16'h0031,16'h003f,16'h0044,-16'h001c,16'h002d,-16'h0072,16'h0015,16'h0037,-16'h002c,-16'h0002,16'h0037,16'h000a,-16'h000f,-16'h0034,-16'h0030,-16'h0021,-16'h0010,16'h0066,16'h0004,16'h005c,16'h002c,16'h0011,16'h0001,-16'h00b6,16'h0037,-16'h0007,16'h0017,-16'h0014,16'h0011,-16'h0020,16'h0014,-16'h0034,-16'h006d,16'h001e,-16'h0033,16'h002a,-16'h0008,16'h0024,16'h0021,-16'h0055,-16'h0029,16'h0024,-16'h0019,16'h0064,16'h002e,-16'h0051,16'h0044,16'h0039,-16'h001a,16'h003f,-16'h0232,16'h002f,-16'h003e,16'h002b,-16'h000e,-16'h0013,-16'h000a,16'h0008,16'h0016,16'h0065,16'h0020,-16'h0036,16'h0012,16'h0016,-16'h0019,16'h0048,16'h0032,16'h0023,16'h0022,-16'h003f,16'h000a,16'h0048,-16'h0067,16'h001e,16'h001f,16'h0009,16'h001e,-16'h0012,-16'h0014,-16'h0051,-16'h0021,16'h0044,16'h0010,16'h0054,16'h0037,16'h0027,16'h0019,-16'h00c5,16'h0039,-16'h0012,16'h0022,-16'h000f,16'h0027,16'h0004,16'h0022,-16'h002a,-16'h0055,16'h0031,-16'h0028,16'h0061,16'h0005,-16'h0008,16'h002e,-16'h0040,16'h0005,16'h0025,16'h002e,16'h003f,16'h0001,-16'h0086,16'h006b,16'h004f,16'h0009,16'h002e,-16'h01f5,16'h0026,-16'h0023,-16'h0006,-16'h0011,16'h0001,16'h003d,16'h0001,16'h0022,16'h0048,16'h0029,-16'h0009,16'h001c,16'h000e,-16'h0044,16'h0043,16'h001e,16'h001c,-16'h00b1,-16'h003f,-16'h0028,16'h0052,-16'h0078,16'h0017,16'h0020,16'h000a,16'h0054,-16'h0027,16'h0039,-16'h0049,-16'h000c,16'h001d,16'h0003,16'h0042,16'h0046,16'h0021,16'h000c,-16'h0123,16'h0055,-16'h0004,16'h000c,-16'h0032,16'h0038,-16'h0002,16'h0007,16'h0001,-16'h0035,16'h0055,16'h0004,16'h004b,16'h0006,-16'h0013,16'h002d,-16'h003c,-16'h000f,16'h0006,-16'h0011,16'h003b,-16'h0005,-16'h007b,16'h0058,16'h0022,-16'h0019,16'h003b,-16'h017c,16'h001f,-16'h0019,16'h000e,-16'h0016,16'h000b,16'h0015,16'h0007,16'h0034,16'h005a,16'h002e,16'h0021,16'h0008,-16'h000c,-16'h0067,16'h005a,16'h000f,-16'h000f,-16'h0229,-16'h0029,16'h001d,16'h005f,-16'h0081,16'h0011,16'h0030,16'h0018,16'h005c,-16'h0006,16'h0035,-16'h004a,-16'h001c,16'h0027,-16'h0009,16'h0042,16'h0065,-16'h000c,16'h001b,-16'h0105,16'h004d,-16'h002c,16'h001c,-16'h0051,16'h0039,16'h000c,-16'h000d,16'h0027,-16'h0002,-16'h0005,16'h002b,16'h005b,16'h0000,-16'h00ad,16'h0038,-16'h0030,-16'h0037,16'h0032,-16'h002a,16'h004f,-16'h0019,-16'h0089,16'h0049,16'h0023,-16'h000e,16'h0025,-16'h0112,16'h0022,-16'h000c,-16'h000d,-16'h0032,16'h002f,16'h0010,16'h0006,16'h0022,16'h0067,16'h001d,16'h002f,-16'h0059,-16'h0015,-16'h00ae,16'h0061,16'h0017,-16'h0037,-16'h026a,-16'h002a,16'h0030,16'h006b,-16'h0085,-16'h0037,16'h003f,16'h005d,16'h0072,-16'h0021,16'h0040,-16'h0005,-16'h0024,-16'h0001,16'h0015,16'h001d,16'h003b,16'h000c,16'h000b,-16'h00c5,16'h001d,-16'h0056,16'h0001,-16'h002f,16'h0065,16'h003c,-16'h000c,16'h0021,-16'h0005,-16'h0024,16'h003f,16'h004d,-16'h0013,-16'h01f5,16'h0006,-16'h003c,16'h002e,16'h002a,-16'h0078,16'h004b,-16'h000d,-16'h0079,16'h0046,16'h0013,-16'h001e,16'h000e,-16'h00d2,16'h0046,16'h000a,16'h0001,-16'h0024,16'h002b,16'h0012,-16'h0002,-16'h0012,16'h004f,16'h0038,-16'h000e,-16'h007e,-16'h0001,-16'h00f0,16'h005e,16'h0005,-16'h0044,-16'h0159,16'h0008,16'h004d,16'h0015,-16'h0070,-16'h0040,16'h0046,16'h003c,16'h0054,16'h0009,16'h002c,16'h003d,-16'h003f,16'h0020,16'h001f,16'h0015,16'h0019,-16'h0007,-16'h0006,-16'h00a3,16'h0029,-16'h0063,-16'h0016,16'h0018,16'h0052,16'h0031,-16'h0008,16'h0018,-16'h000e,-16'h003a,16'h002b,16'h006f,16'h000e,-16'h01bc,16'h001a,-16'h0030,-16'h0011,16'h0032,-16'h0083,16'h0058,16'h000a,-16'h0048,16'h004a,-16'h0008,-16'h001e,-16'h0020,-16'h00b3,16'h0023,16'h0046,16'h001f,-16'h0034,16'h003c,-16'h001c,-16'h0010,16'h000b,16'h004a,16'h0007,16'h0001,-16'h0083,-16'h001e,-16'h00f3,16'h0047,-16'h000d,-16'h0048,-16'h00aa,16'h000d,16'h0027,-16'h00b0,-16'h0037,-16'h0079,16'h0030,-16'h000d,16'h008e,16'h0020,16'h0015,16'h0052,-16'h000f,16'h0031,16'h002a,-16'h0009,16'h0059,-16'h000b,16'h001e,-16'h00a1,16'h0004,-16'h005e,-16'h0035,16'h0058,16'h0033,16'h0034,16'h000f,16'h0049,-16'h0016,-16'h001c,-16'h0017,16'h0064,-16'h0002,-16'h00ea,16'h0031,-16'h002b,-16'h0018,16'h0016,-16'h005c,16'h005e,16'h001b,-16'h002e,16'h0038,-16'h0016,-16'h0012,-16'h005d,-16'h0095,16'h0022,16'h0082,16'h0000,-16'h004c,16'h002a,-16'h0007,-16'h004e,16'h0027,16'h006a,-16'h0018,-16'h0006,-16'h006a,-16'h0033,-16'h00c0,16'h004e,16'h000d,-16'h0036,-16'h005d,16'h003a,16'h0037,-16'h017d,-16'h003c,-16'h0091,16'h0021,-16'h0027,16'h0066,16'h0006,16'h001e,16'h0023,-16'h0030,16'h0022,-16'h0008,16'h0039,16'h0049,16'h0026,16'h001f,-16'h0060,-16'h000c,-16'h004d,-16'h0024,16'h00ba,16'h005e,16'h0055,16'h000b,16'h005b,-16'h0019,-16'h0034,-16'h002a,16'h0047,16'h001e,-16'h0073,16'h0028,-16'h002f,-16'h003c,16'h0006,-16'h0025,16'h0072,16'h0020,-16'h000f,-16'h000c,-16'h0019,-16'h0004,-16'h0062,-16'h0081,-16'h001c,16'h00a8,16'h0000,-16'h005e,16'h0040,16'h0002,-16'h0086,16'h0062,16'h0070,-16'h0026,16'h0011,-16'h007f,-16'h0026,-16'h0078,16'h0046,16'h0012,-16'h003d,16'h0009,16'h0043,16'h002d,-16'h014f,-16'h0021,-16'h006d,16'h0038,-16'h005b,16'h004a,16'h001f,16'h0004,16'h0017,-16'h000b,16'h0034,-16'h0016,16'h003b,16'h0018,16'h0020,16'h0000,-16'h0069,-16'h0012,-16'h001b,-16'h001f,16'h00a5,16'h0063,16'h0036,16'h002f,16'h00a4,16'h0019,-16'h0020,-16'h0018,16'h0042,-16'h0010,-16'h0003,-16'h0025,-16'h003f,-16'h0005,16'h000e,-16'h000f,16'h0058,16'h0008,-16'h003e,-16'h003f,-16'h0008,16'h001a,-16'h0047,-16'h0069,-16'h0023,16'h00b2,16'h0039,-16'h0001,16'h000c,16'h0035,-16'h0052,16'h0065,16'h006f,-16'h0008,16'h0029,-16'h0044,-16'h0014,-16'h0057,16'h003a,-16'h0019,-16'h0008,16'h0024,16'h0053,16'h0049,-16'h00cf,-16'h0003,-16'h0072,16'h0025,-16'h0052,-16'h003d,-16'h0018,16'h001e,16'h001d,16'h0013,16'h0047,16'h000a,16'h00a4,16'h0023,16'h0042,16'h001a,-16'h0055,16'h0000,-16'h0009,-16'h001e,16'h004b,16'h0060,-16'h001b,-16'h0009,16'h0062,16'h000d,-16'h0035,-16'h001c,16'h0026,16'h0010,-16'h0003,-16'h0062,-16'h0034,16'h0026,16'h0068,16'h0028,16'h0013,16'h000b,-16'h0061,16'h0056,16'h0048,-16'h0016,16'h0052,16'h0066,-16'h0002,16'h0077,-16'h0049,16'h0096,-16'h000e,-16'h000f,16'h0027,16'h0013,-16'h001a,-16'h0031,-16'h0062,-16'h003e,16'h002e,16'h005c,-16'h003c,-16'h001c,-16'h005a,16'h003c,-16'h0013,16'h003e,-16'h0027,16'h009f,16'h004d,16'h0019,16'h0000,-16'h001a,-16'h000e,16'h0079,-16'h0029,16'h0014,16'h008a,16'h0019,16'h0016,16'h0013,16'h0002,16'h0021,16'h001c,16'h0004,16'h0030,16'h0060,-16'h002b,16'h0080,16'h0010,16'h001d,16'h003e,-16'h0049,-16'h0018,-16'h0058,-16'h0049,-16'h0052,-16'h0024,16'h0062,16'h0000,16'h0038,16'h0031,16'h0020,16'h002e,16'h0015,-16'h005e,16'h004b,16'h0015,-16'h0014,16'h0041,16'h0067,16'h0003,16'h008c,-16'h0049,16'h0070,-16'h001e,16'h0005,16'h001b,16'h0014,-16'h001b,-16'h0034,-16'h0063,-16'h0055,16'h0010,16'h0061,-16'h0027,-16'h0018,-16'h009f,-16'h0006,-16'h0007,16'h0027,-16'h0003,16'h00c7,16'h007b,16'h0029,16'h000f,-16'h001c,-16'h0021,16'h0037,-16'h0012,-16'h000a,16'h0082,-16'h0005,-16'h0003,-16'h0001,16'h000f,-16'h000a,16'h0015,16'h0002,16'h001e,16'h0019,-16'h001f,16'h0063,16'h0000,16'h0016,16'h005a,-16'h0007,16'h0035,-16'h0041,-16'h0036,-16'h005a,-16'h0027,16'h006f,16'h000b,16'h001d,16'h0027,16'h0011,16'h0027,-16'h000a,-16'h0069,16'h0085,16'h0017,-16'h0015,16'h001f,16'h002c,16'h002c,16'h00bd,-16'h0061,16'h0038,-16'h0002,16'h0037,-16'h0012,16'h002b,-16'h0025,-16'h0054,-16'h0049,-16'h0027,-16'h000b,16'h000b,-16'h001d,16'h0005,-16'h00bc,-16'h0006,-16'h0015,16'h002d,-16'h0001,16'h00d7,16'h0088,16'h0034,-16'h0014,-16'h0035,-16'h000c,16'h0021,-16'h0023,-16'h000c,16'h0076,-16'h000a,16'h0003,-16'h0019,16'h0020,-16'h0039,16'h0028,16'h001b,16'h0011,16'h0027,-16'h0048,16'h001b,-16'h0011,16'h001c,16'h0074,16'h0025,16'h006e,-16'h0005,-16'h0044,-16'h002d,-16'h0011,16'h0036,-16'h0006,16'h002d,16'h0036,16'h001b,16'h003e,-16'h0006,-16'h005e,16'h0048,16'h004b,-16'h0009,16'h0014,16'h0010,16'h005a,16'h0092,-16'h007f,16'h0002,16'h000c,16'h0007,-16'h0009,16'h001d,-16'h0032,-16'h0029,-16'h004e,16'h0000,-16'h0047,16'h0024,16'h0017,16'h001c,-16'h00d0,16'h0019,-16'h002d,16'h000f,-16'h001a,16'h009f,16'h005c,-16'h0007,-16'h0035,-16'h0005,-16'h0015,-16'h0001,-16'h000b,-16'h001f,16'h0091,-16'h004f,-16'h0017,-16'h0015,16'h0017,-16'h0017,16'h0000,16'h0025,16'h0004,16'h0020,-16'h0051,16'h0027,-16'h0017,16'h000e,16'h005e,16'h0058,16'h003b,-16'h001a,-16'h0049,-16'h002a,16'h0010,16'h0024,16'h0000,16'h0044,16'h002a,16'h0030,16'h0044,16'h0002,-16'h0022,16'h0064,16'h0033,16'h0005,-16'h0005,-16'h000d,16'h0059,16'h0067,-16'h004b,-16'h004b,-16'h000a,-16'h0008,-16'h0008,16'h002c,-16'h007b,-16'h0027,-16'h0032,16'h0017,-16'h0065,-16'h0017,16'h0038,16'h003d,-16'h005b,16'h0012,-16'h0039,16'h000b,-16'h000f,16'h0057,16'h0035,16'h0000,-16'h004c,16'h0028,-16'h0018,-16'h004b,-16'h001c,-16'h0038,16'h007d,-16'h005a,16'h000e,-16'h0011,16'h001f,-16'h0021,16'h0009,16'h004e,-16'h003c,16'h0009,-16'h004a,16'h0020,16'h0009,-16'h000c,16'h0054,16'h0044,16'h0011,-16'h0026,-16'h006b,-16'h0027,16'h0003,16'h0011,-16'h0002,16'h0050,-16'h0007,16'h002f,16'h004e,-16'h0021,-16'h0022,16'h0072,16'h004a,16'h0000,16'h0007,-16'h0035,16'h0055,16'h0060,-16'h0042,-16'h0094,16'h0004,16'h0000,-16'h0007,16'h0023,-16'h008d,-16'h0013,-16'h0014,16'h0041,-16'h006a,-16'h0002,16'h003d,16'h0046,-16'h0011,16'h0006,-16'h003b,16'h0006,16'h0040,16'h0061,16'h0030,16'h0022,-16'h002c,16'h0024,-16'h0058,-16'h006a,16'h0001,-16'h000c,16'h0090,-16'h0056,-16'h0017,-16'h0026,16'h0035,-16'h002f,16'h0000,16'h0042,-16'h0038,16'h001b,-16'h004f,16'h0035,-16'h0004,16'h0015,16'h005f,16'h005f,-16'h0001,-16'h001b,-16'h009f,-16'h0015,16'h000f,16'h004e,-16'h0027,16'h0034,-16'h0016,16'h0027,16'h004e,-16'h003c,16'h0002,16'h0070,16'h0049,16'h0005,-16'h0013,-16'h001f,16'h0067,16'h0028,-16'h0025,-16'h00c2,16'h001d,-16'h0007,-16'h0024,16'h0016,-16'h008b,-16'h002b,16'h0000,16'h004c,-16'h0051,16'h0012,16'h0068,16'h0035,-16'h002c,-16'h0015,-16'h0026,-16'h0026,16'h0038,16'h0069,16'h0020,16'h0024,-16'h0010,16'h0041,-16'h008b,-16'h005b,16'h0033,-16'h001e,16'h008a,16'h0001,-16'h0032,-16'h0026,16'h0013,-16'h000f,16'h0000,16'h001b,-16'h000b,16'h000e,-16'h0002,16'h0036,-16'h000a,16'h0012,16'h000f,16'h0015,-16'h001b,-16'h0042,-16'h009f,-16'h002f,-16'h0019,16'h0051,-16'h000c,16'h0033,-16'h0002,16'h0012,16'h004b,-16'h0050,-16'h0007,16'h0080,16'h0054,16'h0001,-16'h000f,-16'h0035,16'h007e,16'h0015,16'h0010,-16'h00c1,16'h002b,16'h0017,16'h0006,16'h0032,-16'h005d,-16'h0030,16'h0002,16'h003d,-16'h0021,16'h0024,16'h005e,16'h0025,-16'h003c,16'h0003,-16'h0028,-16'h004a,16'h0029,16'h0063,16'h0017,16'h001e,16'h0018,-16'h000c,-16'h0051,-16'h0029,16'h0050,-16'h003e,16'h00a4,16'h0032,-16'h0051,-16'h0021,16'h000f,16'h0013,-16'h0004,16'h0022,-16'h001e,16'h0020,16'h0011,16'h002d,-16'h0023,16'h0038,16'h0000,16'h000d,-16'h004d,-16'h0015,-16'h00c4,-16'h0017,-16'h0006,16'h0030,-16'h004b,16'h0026,-16'h0006,16'h001b,16'h005b,-16'h00b0,-16'h000a,16'h0080,16'h004e,-16'h000a,16'h0002,-16'h007f,16'h0077,16'h0019,16'h002a,-16'h00d6,16'h0014,16'h0019,-16'h000b,16'h0025,-16'h003b,-16'h0033,16'h000c,16'h0006,16'h0000,16'h0025,16'h0042,16'h0004,-16'h0049,-16'h0010,-16'h0044,-16'h0043,16'h001e,16'h0067,16'h003d,16'h0003,16'h0030,-16'h0044,-16'h001c,16'h0007,16'h0039,-16'h0023,16'h0097,-16'h000c,-16'h0056,-16'h0030,16'h0004,16'h000b,16'h0007,16'h0020,-16'h0035,16'h0021,16'h0026,-16'h0016,-16'h0016,16'h001d,-16'h000a,16'h000e,-16'h0032,16'h000b,-16'h00e8,-16'h0005,-16'h000c,16'h004d,-16'h0022,16'h0052,-16'h0028,-16'h0003,16'h0057,-16'h00b1,-16'h001b,16'h0081,16'h0068,-16'h0008,-16'h0017,-16'h009a,16'h008d,16'h001f,16'h0037,-16'h00f1,-16'h0005,16'h0033,-16'h0001,-16'h0012,-16'h0036,-16'h0025,16'h0007,16'h0012,-16'h0027,16'h002d,16'h005b,-16'h0055,-16'h0009,-16'h0018,-16'h0024,-16'h000c,16'h0028,16'h005d,16'h0025,16'h0012,16'h0024,-16'h0052,-16'h000e,-16'h0005,-16'h0037,-16'h0006,16'h005f,16'h0004,-16'h0042,-16'h004c,16'h0020,16'h0015,-16'h0004,16'h0036,-16'h000b,16'h001f,16'h0018,16'h000c,-16'h0028,16'h0025,-16'h003b,16'h0024,-16'h0011,16'h0002,-16'h00fb,16'h0018,16'h000a,16'h0034,-16'h0019,16'h0060,-16'h004a,-16'h0028,16'h0084,-16'h00a3,-16'h0006,16'h008e,16'h0048,-16'h0026,-16'h0009,-16'h00d9,16'h008f,16'h000e,16'h001b,-16'h0150,-16'h002e,16'h0034,-16'h0008,-16'h001b,-16'h002c,-16'h000f,-16'h0016,16'h0002,-16'h0016,-16'h0001,16'h005c,-16'h005c,-16'h0001,16'h0001,-16'h005c,16'h0012,16'h001b,16'h006f,-16'h0020,16'h0036,16'h001c,-16'h000c,16'h0008,16'h0004,-16'h00a3,-16'h0044,16'h005f,16'h0002,-16'h003d,-16'h0050,-16'h0008,16'h001d,-16'h0006,16'h0023,16'h0006,16'h001d,-16'h000c,-16'h0005,-16'h004a,16'h0038,-16'h0031,16'h000a,16'h002a,16'h0028,-16'h00dd,-16'h0003,16'h003b,16'h0019,-16'h001c,16'h0026,-16'h003f,-16'h000e,16'h0037,-16'h009e,-16'h0016,16'h009c,16'h0028,-16'h0028,16'h0017,-16'h0104,16'h00a7,16'h0000,16'h004d,-16'h015c,-16'h0011,16'h000d,16'h0019,16'h0035,-16'h0017,-16'h0009,-16'h0029,16'h002c,-16'h0018,16'h000d,16'h0065,-16'h0023,-16'h0014,16'h001f,-16'h005f,16'h003c,16'h000d,16'h0068,-16'h0076,16'h0037,16'h0034,16'h001b,-16'h003c,16'h000a,-16'h0079,-16'h0046,16'h0067,-16'h0009,-16'h000b,-16'h0067,-16'h0017,16'h0046,-16'h0029,16'h001d,-16'h0009,16'h001e,-16'h0015,16'h0018,-16'h0042,16'h0013,-16'h0019,-16'h0002,16'h0019,-16'h000f,-16'h00d8,-16'h0008,16'h003d,16'h0026,-16'h0039,-16'h0006,-16'h0059,-16'h000b,16'h001e,-16'h0099,16'h0007,16'h00a6,16'h002f,-16'h001a,16'h002e,-16'h0143,16'h0080,-16'h0039,16'h003e,-16'h019c,16'h0012,16'h0027,16'h0011,16'h003c,16'h0005,-16'h0025,16'h000e,16'h0012,16'h0007,-16'h0001,16'h0070,-16'h003b,-16'h002a,16'h0007,-16'h0060,16'h003f,-16'h0011,16'h002f,-16'h0093,16'h0012,16'h0016,16'h0000,-16'h0031,-16'h0031,-16'h004d,-16'h0028,16'h0044,-16'h000e,-16'h0003,-16'h009e,-16'h0039,16'h0037,-16'h0043,16'h001a,-16'h0008,16'h002a,-16'h0028,16'h0020,-16'h003e,16'h001a,-16'h001b,-16'h0002,16'h0034,16'h000b,-16'h0090,16'h0014,16'h0029,-16'h000a,-16'h0014,16'h000a,-16'h004f,16'h0021,16'h0015,-16'h00ac,-16'h001d,16'h00a3,16'h002c,-16'h0022,16'h0054,-16'h0151,16'h0079,-16'h000f,16'h0039,-16'h01e0,16'h000e,16'h001f,-16'h0004,16'h002a,16'h0028,-16'h0028,16'h0002,16'h002b,16'h0023,-16'h000c,16'h0051,-16'h0018,-16'h0052,16'h0009,-16'h0067,16'h0047,-16'h0027,-16'h0013,-16'h006c,16'h0013,16'h0004,-16'h001a,16'h0003,-16'h0047,-16'h0021,-16'h000f,16'h002d,-16'h0026,-16'h0031,-16'h0055,-16'h002c,16'h0021,-16'h0040,16'h002b,-16'h0014,16'h0020,-16'h003b,16'h0033,-16'h003f,-16'h0002,-16'h001c,-16'h0030,16'h0000,-16'h0013,-16'h0031,16'h001b,16'h0038,-16'h0008,-16'h002d,-16'h001e,-16'h0033,16'h001f,16'h002a,-16'h0098,-16'h0008,16'h0082,16'h0029,-16'h002d,16'h0026,-16'h0140,16'h006b,16'h0008,16'h0064,-16'h01fc,-16'h001a,-16'h0007,-16'h0004,16'h000f,16'h002f,-16'h0008,16'h003b,16'h0018,16'h0030,16'h001e,16'h0065,16'h0029,-16'h0064,16'h0026,-16'h0071,16'h0050,-16'h0014,-16'h001d,-16'h0043,16'h000d,16'h0022,-16'h0027,16'h001c,-16'h0026,16'h003d,-16'h0022,16'h0018,-16'h002d,-16'h0020,-16'h002c,-16'h0013,16'h0031,-16'h003c,16'h0045,-16'h0007,16'h0041,-16'h0029,16'h0045,-16'h0032,-16'h0006,-16'h0013,-16'h0007,-16'h0067,-16'h0009,16'h0029,16'h0005,16'h0033,-16'h0009,-16'h0048,-16'h0016,-16'h001a,16'h0024,16'h0033,-16'h008a,-16'h0003,16'h007e,16'h0026,-16'h0002,16'h0003,-16'h0169,16'h006a,-16'h0016,16'h0041,-16'h01e2,-16'h0037,-16'h003a,-16'h0012,16'h0021,16'h0025,-16'h0007,16'h0026,16'h0015,16'h0004,16'h0009,16'h0072,16'h002c,-16'h0026,16'h0054,-16'h00b0,16'h0017,-16'h0032,-16'h0012,16'h0000,16'h0007,16'h0017,-16'h0039,16'h0038,-16'h002e,16'h003f,16'h0006,16'h0030,-16'h002c,-16'h004d,16'h002d,-16'h0033,16'h004a,-16'h001a,16'h002f,-16'h0019,16'h0050,-16'h0026,16'h0054,-16'h0016,-16'h000b,-16'h0013,-16'h0006,-16'h009a,-16'h002f,16'h000d,16'h0013,16'h0009,16'h0008,-16'h004e,-16'h0007,16'h0003,16'h0006,16'h0040,-16'h0089,-16'h0018,16'h0068,16'h003e,-16'h0014,-16'h000e,-16'h017a,16'h004c,-16'h000a,16'h0036,-16'h01ba,-16'h0030,-16'h0020,-16'h0034,-16'h000d,16'h0047,16'h0013,16'h001c,16'h002b,-16'h001b,16'h000e,16'h0058,16'h001b,16'h0003,16'h0060,-16'h00a4,-16'h0061,-16'h0032,-16'h0008,16'h0006,16'h0036,16'h0009,-16'h005b,16'h001c,-16'h003e,16'h0040,16'h000a,16'h0042,-16'h0025,-16'h001d,16'h005e,-16'h000c,16'h0048,-16'h0049,16'h003f,16'h0006,16'h0043,-16'h0017,16'h002e,-16'h0018,16'h000c,-16'h0049,16'h001f,-16'h008a,-16'h0053,-16'h000d,16'h0023,16'h0024,16'h0008,-16'h002b,16'h000c,16'h0002,-16'h0025,16'h0059,-16'h007f,-16'h001a,16'h0042,16'h0044,-16'h0024,-16'h0007,-16'h019a,16'h002d,-16'h0012,16'h001e,-16'h018d,-16'h000e,-16'h000f,-16'h0028,16'h0007,16'h0034,16'h0012,16'h0010,16'h0023,-16'h000f,16'h0011,16'h0054,16'h0040,-16'h0020,16'h0064,-16'h0086,-16'h000c,16'h000e,-16'h0033,16'h0025,16'h0021,-16'h0014,-16'h0023,16'h0011,-16'h0044,-16'h0001,16'h0021,16'h0050,-16'h0015,16'h0025,16'h0075,-16'h0015,16'h0006,-16'h00a1,16'h0019,-16'h0025,16'h0043,-16'h001c,16'h0034,-16'h0006,16'h000e,-16'h0040,-16'h0011,-16'h001b,-16'h006a,16'h001e,-16'h0004,-16'h0008,16'h0028,-16'h001b,-16'h0015,-16'h0003,-16'h001d,16'h004c,-16'h003f,-16'h0031,16'h006c,16'h003b,-16'h001f,16'h0019,-16'h01b7,16'h000a,-16'h002a,16'h0024,-16'h0153,16'h0001,16'h0000,-16'h001d,16'h0018,16'h0059,16'h002d,-16'h000c,16'h0025,16'h0002,-16'h0017,16'h0060,16'h0029,16'h0001,16'h0043,-16'h00ae,-16'h0007,16'h0033,-16'h0077,16'h001a,16'h0027,-16'h000e,16'h0000,-16'h0026,-16'h001e,-16'h0030,16'h0000,16'h0026,-16'h000f,16'h0056,16'h0061,-16'h000f,16'h0002,-16'h0111,16'h0034,-16'h0029,16'h0017,-16'h0030,16'h0027,16'h0002,-16'h000a,-16'h003b,-16'h0031,16'h0028,-16'h0040,16'h0031,16'h0036,16'h0021,-16'h0012,-16'h0037,16'h0018,16'h0016,16'h0014,16'h0056,-16'h000c,-16'h005d,16'h005a,16'h004a,-16'h000a,16'h002d,-16'h019e,16'h0027,-16'h0046,16'h0024,-16'h012a,16'h0004,16'h0017,-16'h000a,16'h0028,16'h004a,16'h0020,-16'h002c,16'h003d,16'h0000,-16'h004a,16'h0037,16'h001c,16'h003a,16'h0037,-16'h00d0,16'h0019,16'h003f,-16'h00ab,16'h0022,16'h0019,16'h000a,16'h001f,-16'h001b,-16'h0003,-16'h0081,-16'h0016,16'h0037,-16'h0012,16'h0045,16'h0054,-16'h0014,16'h0006,-16'h0131,16'h0023,-16'h0030,-16'h0011,-16'h0043,16'h0031,16'h0012,16'h0016,-16'h0013,-16'h0022,16'h0047,-16'h0038,16'h0048,16'h004c,-16'h002e,-16'h0002,-16'h0012,16'h0014,16'h001b,16'h0013,16'h0063,-16'h001c,-16'h0069,16'h005d,16'h004a,-16'h0004,16'h002e,-16'h0156,16'h0022,-16'h005b,16'h0019,-16'h010e,16'h000c,16'h0049,-16'h001a,16'h0042,16'h0056,16'h0019,-16'h0018,16'h0053,-16'h0012,-16'h0052,16'h0034,16'h0001,16'h0029,-16'h00bd,-16'h00ba,16'h0001,16'h0069,-16'h00d1,-16'h000b,16'h0025,16'h0023,16'h0079,-16'h001b,16'h0037,-16'h0067,-16'h0023,16'h0009,16'h0014,16'h0046,16'h004c,-16'h0026,16'h0004,-16'h0151,16'h001c,-16'h0016,-16'h0010,-16'h0055,16'h002f,16'h003b,-16'h0015,16'h0017,-16'h0014,16'h0038,-16'h0001,16'h0061,16'h002c,-16'h006b,16'h0010,16'h0007,-16'h0017,16'h0040,-16'h0018,16'h0042,-16'h0006,-16'h0079,16'h0053,16'h001c,-16'h0021,16'h002d,-16'h00f8,16'h004b,-16'h0024,16'h0005,-16'h00fc,16'h0025,16'h000f,16'h0006,16'h0030,16'h004d,16'h0005,16'h001b,16'h0042,-16'h0024,-16'h008d,16'h001f,-16'h0022,-16'h000e,-16'h0206,-16'h00c8,16'h000e,16'h004e,-16'h00aa,-16'h0046,16'h0002,16'h003b,16'h007c,-16'h000f,16'h0043,-16'h0028,-16'h000d,16'h0008,16'h0003,16'h002b,16'h0047,-16'h0061,-16'h000d,-16'h00e1,16'h0003,-16'h0042,16'h0019,-16'h004e,16'h003d,16'h0061,-16'h0011,16'h0023,16'h0001,16'h0006,16'h001f,16'h0078,16'h0006,-16'h0112,16'h002b,-16'h0009,-16'h0016,16'h0024,-16'h006a,16'h0063,16'h000d,-16'h007a,16'h0049,16'h001f,-16'h0033,16'h0019,-16'h00ae,16'h0035,-16'h0012,16'h001f,-16'h00ec,16'h000b,16'h003b,-16'h000e,16'h0009,16'h007b,16'h0009,16'h0003,-16'h000b,-16'h0023,-16'h00d3,16'h005e,-16'h002c,-16'h002d,-16'h022d,-16'h00ba,16'h002c,16'h003b,-16'h007e,-16'h0057,16'h0013,16'h006e,16'h007e,-16'h000a,16'h0049,16'h0029,-16'h0015,16'h002b,16'h002b,16'h005a,16'h0036,-16'h001d,-16'h0006,-16'h009b,-16'h0006,-16'h0058,16'h0001,-16'h002e,16'h0071,16'h004e,16'h0001,-16'h0017,16'h0000,-16'h0036,16'h0026,16'h006f,16'h002f,-16'h01b2,16'h0021,16'h0008,-16'h0009,16'h004a,-16'h00a0,16'h0040,16'h0036,-16'h0050,16'h004d,-16'h0004,-16'h001c,-16'h000f,-16'h0093,16'h0044,16'h0008,16'h001a,-16'h00c9,16'h0027,16'h0025,-16'h0041,-16'h003f,16'h0059,-16'h0012,-16'h0028,-16'h0034,-16'h0007,-16'h00d5,16'h006b,-16'h0027,-16'h0048,-16'h0136,-16'h00b1,16'h0030,16'h0000,-16'h0059,-16'h0068,16'h0043,16'h0056,16'h009d,16'h000c,16'h0044,16'h003f,-16'h000f,16'h0032,16'h002b,16'h002c,16'h0037,-16'h0013,16'h000b,-16'h0072,16'h0001,-16'h0068,-16'h0015,16'h001a,16'h0059,16'h003f,-16'h0022,16'h0006,-16'h000c,-16'h0047,16'h002b,16'h0066,-16'h0004,-16'h013e,16'h0037,16'h0004,-16'h001c,-16'h0008,-16'h008a,16'h005b,16'h001c,-16'h001a,16'h004d,16'h0001,-16'h0016,-16'h002d,-16'h006d,16'h001b,16'h005b,16'h0023,-16'h00ce,16'h0013,16'h0036,-16'h0012,-16'h0015,16'h0064,16'h0004,-16'h0001,-16'h0027,-16'h0016,-16'h00d0,16'h0063,16'h0004,-16'h005c,-16'h009f,-16'h0079,16'h002e,-16'h00b2,-16'h0037,-16'h0060,16'h0029,-16'h0008,16'h0072,16'h001d,16'h002b,16'h005f,-16'h0017,16'h0043,-16'h000e,16'h0019,16'h0016,16'h001b,16'h0001,-16'h0077,16'h0003,-16'h005f,-16'h0050,16'h0083,16'h005b,16'h003c,16'h000d,16'h0011,16'h0003,-16'h005e,-16'h000a,16'h0082,-16'h0016,-16'h0097,16'h003f,-16'h000d,-16'h004b,-16'h0005,-16'h004a,16'h0063,16'h003f,-16'h001d,16'h003c,-16'h000a,-16'h0013,-16'h005b,-16'h007f,16'h0004,16'h009b,16'h0005,-16'h00b8,16'h0019,16'h0027,-16'h0054,16'h002d,16'h0061,-16'h000a,16'h0013,-16'h005a,16'h0003,-16'h00aa,16'h0054,-16'h0017,-16'h0053,-16'h004b,-16'h0063,16'h004e,-16'h0138,-16'h0024,-16'h0067,16'h0013,-16'h0016,16'h0076,16'h0014,16'h0001,16'h0047,-16'h0013,16'h0036,-16'h001c,16'h0055,16'h0034,16'h0023,16'h0011,-16'h0062,16'h0000,-16'h0038,-16'h0038,16'h008f,16'h0068,16'h0032,16'h0016,16'h0034,-16'h0004,-16'h0040,-16'h0026,16'h0051,-16'h0015,-16'h005a,16'h0003,-16'h0014,-16'h0033,-16'h0013,-16'h002c,16'h005b,16'h000e,-16'h0013,-16'h0005,-16'h000b,16'h0006,-16'h006a,-16'h0058,-16'h0032,16'h009e,16'h0014,-16'h008a,16'h003c,16'h000a,-16'h0045,16'h003b,16'h0079,16'h000c,16'h0020,-16'h005d,-16'h000d,-16'h005b,16'h0051,-16'h0001,-16'h004e,-16'h0003,-16'h0025,16'h0062,-16'h00fc,16'h0001,-16'h0080,16'h0024,-16'h0038,16'h0018,16'h0018,-16'h0009,16'h0037,-16'h001e,16'h002e,-16'h000c,16'h006f,-16'h0006,16'h0023,16'h0027,-16'h003a,16'h0016,-16'h0014,-16'h0021,16'h006d,16'h0050,16'h0007,-16'h0014,16'h0033,16'h002b,-16'h000e,-16'h001f,16'h004b,-16'h0011,16'h0000,-16'h0023,16'h0003,16'h0008,-16'h0028,-16'h0027,16'h004c,16'h0002,-16'h0061,-16'h000d,-16'h0009,16'h0041,-16'h0045,-16'h0068,-16'h0031,16'h00a1,16'h0038,-16'h0033,-16'h0011,16'h0018,-16'h0042,16'h0058,16'h0092,16'h000b,16'h0023,-16'h002b,16'h001c,-16'h0035,16'h0054,-16'h0010,-16'h002a,16'h0014,16'h0002,16'h004d,-16'h009f,-16'h000f,-16'h006c,16'h0016,-16'h000a,-16'h0037,16'h0007,-16'h0012,16'h004a,-16'h0001,16'h0043,-16'h000e,16'h00ae,-16'h0018,16'h001a,16'h000e,-16'h0047,16'h000b,-16'h000a,-16'h0013,16'h003f,16'h0063,-16'h0020,-16'h004b,16'h003b,16'h002c,-16'h003b,-16'h0036,16'h004b,16'h0025,-16'h0008,-16'h0049,-16'h0030,16'h0042,16'h0045,16'h000f,16'h0032,16'h000d,-16'h0046,16'h0045,16'h003b,-16'h001b,16'h005a,16'h0050,16'h0014,16'h0061,-16'h003d,16'h000e,-16'h0025,-16'h0014,16'h004f,-16'h0011,-16'h0016,-16'h002e,-16'h0033,-16'h0036,16'h002a,16'h0046,-16'h002d,-16'h0003,-16'h0056,16'h001f,-16'h0008,16'h0039,-16'h0028,16'h0078,16'h0035,-16'h000e,16'h0015,16'h0001,-16'h0016,16'h005e,-16'h0018,16'h0006,16'h0070,-16'h0016,-16'h0004,16'h0010,-16'h0008,16'h0002,16'h002c,-16'h000b,16'h0020,16'h0055,-16'h0017,16'h0068,16'h0011,16'h0019,16'h0028,-16'h0040,-16'h0027,-16'h0055,-16'h0011,-16'h0033,-16'h0027,16'h002f,-16'h0018,16'h0033,16'h002e,-16'h0001,16'h0025,-16'h000a,-16'h005e,16'h0053,16'h002b,-16'h0021,16'h0045,16'h004e,16'h001c,16'h0079,-16'h0033,16'h0015,16'h0005,16'h0019,16'h003f,16'h0018,16'h000c,-16'h001f,-16'h004f,-16'h005d,16'h002e,16'h0037,-16'h001c,-16'h0001,-16'h005f,16'h0010,16'h0006,16'h0027,-16'h001d,16'h0080,16'h0065,16'h0005,-16'h0003,16'h001a,-16'h0008,16'h0039,-16'h001e,16'h000e,16'h0065,-16'h0005,-16'h0009,-16'h0005,-16'h000d,-16'h0003,16'h000b,16'h0002,16'h0039,16'h002d,-16'h003c,16'h0042,-16'h000b,16'h0010,16'h0050,-16'h0028,-16'h0010,-16'h005f,-16'h0028,-16'h0052,16'h0000,16'h0032,16'h000f,16'h0029,16'h0046,16'h000c,16'h0021,16'h000b,-16'h004f,16'h0080,16'h001d,-16'h0026,16'h0043,16'h0041,16'h0018,16'h00a1,-16'h0068,16'h0037,-16'h0008,16'h0011,16'h0022,16'h0006,-16'h001b,-16'h001d,-16'h0052,-16'h0039,16'h001b,16'h002c,-16'h000f,16'h0012,-16'h0090,16'h001b,-16'h0018,16'h0028,16'h001f,16'h00ad,16'h0071,16'h001f,-16'h0021,16'h000c,-16'h0017,16'h003c,-16'h0026,-16'h0024,16'h0063,-16'h0021,-16'h0001,-16'h003b,16'h000c,16'h0009,16'h0023,16'h0000,16'h0027,16'h002e,-16'h0031,16'h0025,-16'h000c,-16'h0008,16'h0072,16'h0002,16'h001a,-16'h0031,-16'h002a,-16'h0024,16'h0004,16'h0026,16'h0007,16'h0010,16'h0055,16'h000c,16'h001c,-16'h0011,-16'h004c,16'h006f,16'h0008,-16'h001c,16'h002c,16'h0003,16'h0023,16'h008e,-16'h0065,-16'h000a,16'h0006,16'h0000,16'h0000,16'h0004,-16'h0021,-16'h001f,-16'h0050,-16'h0021,-16'h000a,16'h0009,16'h0001,-16'h0006,-16'h0066,16'h000f,-16'h0010,16'h0020,16'h000d,16'h00d0,16'h0085,-16'h0007,-16'h002c,16'h0028,-16'h001a,16'h002d,-16'h000d,-16'h0023,16'h0063,-16'h0054,-16'h0013,-16'h004a,16'h0002,-16'h0044,16'h0016,16'h0002,16'h0014,16'h0028,-16'h0058,16'h0025,-16'h0014,-16'h000d,16'h004c,16'h000d,16'h002b,-16'h0043,-16'h0048,-16'h0030,16'h000d,16'h0012,-16'h0010,16'h0030,16'h003d,16'h000f,16'h0030,-16'h001f,-16'h0025,16'h006d,16'h0020,-16'h0009,16'h003b,-16'h0027,16'h0032,16'h008f,-16'h004a,-16'h0076,-16'h0003,-16'h000d,16'h0005,16'h0012,-16'h005e,-16'h0015,-16'h004b,16'h0016,-16'h0049,16'h0010,16'h001e,16'h000e,-16'h0061,16'h0000,16'h0000,-16'h0005,16'h001e,16'h007d,16'h003e,16'h000f,-16'h0062,16'h0053,-16'h0022,-16'h0012,-16'h0019,-16'h0037,16'h0082,-16'h0060,-16'h0027,-16'h004d,16'h000f,-16'h003b,16'h0021,16'h0000,-16'h0027,16'h001c,-16'h005b,16'h0025,-16'h0012,16'h0006,16'h0030,16'h0001,16'h0011,-16'h0049,-16'h0072,-16'h000e,16'h0002,16'h0028,-16'h0005,16'h003b,16'h001a,16'h0029,16'h0058,-16'h001c,16'h001b,16'h0069,16'h001f,16'h000e,16'h0012,-16'h0053,16'h0032,16'h007e,-16'h002c,-16'h00ca,16'h001b,16'h0005,16'h0002,16'h0025,-16'h0081,16'h0013,-16'h001e,16'h003c,-16'h0059,-16'h0002,16'h0015,16'h004c,-16'h0017,-16'h0003,16'h0000,-16'h001f,16'h003e,16'h008c,16'h003b,16'h000a,-16'h0035,16'h006f,-16'h004a,-16'h0041,16'h000a,-16'h0025,16'h0086,-16'h0056,-16'h0029,-16'h003b,16'h0019,-16'h0038,16'h0019,16'h0018,-16'h003f,16'h0010,-16'h0036,16'h002f,-16'h0022,-16'h0011,16'h001e,16'h0006,16'h0023,-16'h003a,-16'h009d,16'h0005,-16'h0011,16'h0035,16'h0015,16'h002f,16'h0028,16'h000c,16'h0040,-16'h0069,16'h0031,16'h0066,16'h001d,-16'h000c,-16'h0003,-16'h0071,16'h0034,16'h004d,-16'h0031,-16'h00d9,16'h0015,16'h0010,16'h0004,16'h0005,-16'h007a,-16'h000c,16'h0006,16'h005b,-16'h002b,16'h002d,16'h0030,16'h0049,-16'h003e,-16'h0011,-16'h000c,-16'h0030,16'h0046,16'h0049,-16'h0014,16'h0004,-16'h0024,16'h006a,-16'h007a,-16'h0032,16'h0036,-16'h0047,16'h0094,16'h0018,-16'h0020,-16'h0047,16'h0015,-16'h0022,16'h0002,16'h001e,-16'h0041,16'h0005,16'h0017,16'h0049,16'h0000,-16'h000d,-16'h000b,16'h0018,16'h002f,-16'h0048,-16'h00f6,-16'h0015,16'h0004,16'h0053,-16'h0007,16'h002b,16'h0001,16'h0004,16'h0069,-16'h00ad,16'h0036,16'h007f,16'h004f,16'h0014,-16'h000c,-16'h00ad,16'h004f,16'h0032,-16'h0002,-16'h0125,16'h000c,16'h0036,-16'h0014,-16'h0009,-16'h0074,-16'h0017,-16'h002a,16'h0053,-16'h0030,16'h0016,16'h0046,16'h0022,-16'h0030,-16'h0009,-16'h000b,-16'h0064,16'h0044,16'h0059,-16'h001a,16'h002a,-16'h0002,16'h0043,-16'h0052,-16'h0043,16'h0034,-16'h004d,16'h007e,16'h001b,-16'h004d,-16'h0039,-16'h000c,16'h0015,-16'h0005,-16'h0005,-16'h0039,16'h0028,16'h0016,16'h0039,-16'h0003,16'h0009,-16'h0037,16'h0004,16'h0001,-16'h0044,-16'h011e,-16'h0007,16'h0000,16'h004d,-16'h001e,16'h0049,-16'h000a,16'h000e,16'h004f,-16'h00f2,16'h0018,16'h0049,16'h0055,16'h0002,-16'h0022,-16'h00e8,16'h005d,16'h0039,16'h0020,-16'h0193,16'h001b,16'h0021,-16'h0001,-16'h0009,-16'h0082,-16'h0021,-16'h0003,16'h0033,16'h0000,16'h0033,16'h003a,-16'h0002,-16'h0016,-16'h0013,-16'h0029,-16'h0047,16'h0015,16'h0041,-16'h0004,-16'h0005,16'h0006,-16'h001f,-16'h0014,-16'h0003,-16'h0002,-16'h001e,16'h008e,16'h0037,-16'h0054,-16'h0020,-16'h0008,16'h0013,16'h0027,16'h0010,-16'h0021,16'h0011,16'h0020,16'h0017,-16'h0012,16'h0018,-16'h003c,-16'h0019,16'h0015,-16'h001f,-16'h0111,16'h0031,16'h0040,16'h0036,-16'h0036,16'h002d,-16'h0019,16'h000b,16'h0058,-16'h0128,16'h0027,16'h0054,16'h0087,-16'h0007,-16'h0021,-16'h0107,16'h006e,16'h001f,16'h0026,-16'h0217,16'h0023,16'h0031,16'h001b,-16'h005d,-16'h0072,-16'h0021,16'h001d,16'h0000,16'h0003,16'h0036,16'h003c,-16'h0079,16'h0005,-16'h0004,-16'h001c,-16'h002d,16'h0014,16'h003c,16'h000c,16'h000b,16'h001b,-16'h0035,16'h0036,16'h0000,-16'h0037,-16'h001f,16'h0067,16'h001b,-16'h0014,-16'h003e,-16'h0006,16'h001e,16'h0011,16'h002b,-16'h000c,-16'h0005,16'h0034,16'h002e,-16'h000c,16'h0017,-16'h0045,-16'h000a,16'h000e,-16'h0016,-16'h00f4,16'h001d,16'h0020,16'h0028,-16'h0039,16'h002e,-16'h0036,-16'h0017,16'h0059,-16'h0109,16'h003c,16'h003a,16'h004e,-16'h0002,-16'h002b,-16'h00e3,16'h0069,16'h0029,16'h0020,-16'h0248,-16'h0016,16'h0035,16'h0015,-16'h0025,-16'h0082,16'h0013,-16'h003d,16'h001f,16'h0006,16'h0015,16'h0039,-16'h005d,16'h002f,16'h0014,-16'h002c,16'h001a,-16'h0009,16'h0002,-16'h0021,16'h0034,16'h002b,-16'h000e,16'h0009,-16'h0004,-16'h0070,-16'h0018,16'h005b,-16'h0005,-16'h0028,-16'h005b,16'h0010,16'h0000,16'h0010,16'h002f,16'h000b,-16'h0009,16'h002a,16'h001f,-16'h0026,16'h0035,-16'h001d,16'h0000,16'h0037,-16'h0032,-16'h0103,16'h002d,16'h003b,16'h0025,-16'h002d,16'h0035,-16'h001a,-16'h003d,16'h004e,-16'h00fd,16'h0042,16'h004c,16'h0048,-16'h0010,16'h0017,-16'h0102,16'h0078,-16'h0019,16'h0033,-16'h028f,-16'h000f,16'h001a,16'h0023,16'h0024,-16'h0064,16'h0016,-16'h002f,16'h0025,-16'h0001,-16'h000c,16'h0048,-16'h0028,16'h0031,16'h0011,-16'h0043,16'h0027,-16'h0021,16'h000d,-16'h005c,16'h002f,16'h0023,16'h0007,-16'h0038,-16'h0004,-16'h004a,-16'h0012,16'h0064,16'h001d,16'h0014,-16'h004e,-16'h0002,16'h0024,16'h0006,16'h0032,-16'h0016,-16'h0009,-16'h0039,16'h001b,-16'h002d,16'h0038,-16'h0014,-16'h001e,16'h0031,-16'h0029,-16'h0103,16'h0011,16'h0023,16'h0006,-16'h0030,-16'h001e,-16'h0009,-16'h0028,16'h0030,-16'h00ed,16'h0033,16'h004b,16'h0032,-16'h001f,16'h0059,-16'h00cc,16'h006d,-16'h002f,16'h0049,-16'h0272,-16'h0001,16'h0004,16'h001e,16'h0048,-16'h0054,16'h0018,16'h001d,16'h001b,16'h0002,16'h0001,16'h0023,-16'h0021,-16'h0005,16'h0003,-16'h005f,16'h004f,-16'h002a,-16'h0005,-16'h006d,16'h0032,-16'h0011,-16'h0005,-16'h003e,-16'h002a,-16'h0041,-16'h0014,16'h007e,16'h0002,16'h0012,-16'h0067,-16'h0026,16'h002a,16'h000a,16'h0018,-16'h001c,16'h0012,-16'h002e,16'h0027,-16'h002a,16'h0024,-16'h0031,-16'h0016,16'h0015,-16'h0041,-16'h0128,16'h0013,16'h0040,-16'h0001,-16'h0016,-16'h002d,-16'h0021,-16'h000f,16'h003e,-16'h00da,-16'h0003,16'h0071,16'h0035,-16'h001b,16'h0044,-16'h00a2,16'h004f,-16'h000c,16'h0046,-16'h0222,-16'h000a,16'h0009,16'h0018,16'h002f,-16'h003c,16'h000a,16'h0041,16'h0017,16'h002b,16'h0001,16'h0040,16'h0003,-16'h0042,16'h0002,-16'h004a,16'h0040,-16'h0027,-16'h0027,-16'h0036,16'h0026,-16'h0002,-16'h000b,16'h0000,-16'h005a,-16'h002c,16'h000d,16'h005a,-16'h0015,-16'h0005,-16'h0051,-16'h001c,16'h001b,-16'h0045,16'h0012,-16'h0013,16'h0028,-16'h0016,16'h0047,-16'h0025,16'h002e,-16'h002a,-16'h000a,-16'h0001,-16'h0024,-16'h00d2,-16'h000e,16'h0014,-16'h000f,-16'h0016,-16'h000f,16'h0005,16'h0022,16'h003b,-16'h00bb,16'h0000,16'h0062,16'h0045,-16'h002e,16'h0039,-16'h0094,16'h0058,16'h000b,16'h003e,-16'h021f,-16'h002b,-16'h001a,-16'h0007,16'h001d,-16'h0020,16'h0005,16'h001a,16'h001d,16'h002b,-16'h0023,16'h004b,16'h0031,-16'h002d,16'h0020,-16'h0054,16'h004b,-16'h002d,-16'h0042,-16'h0004,16'h0023,16'h000d,-16'h0015,16'h002d,-16'h0030,16'h0042,16'h0000,16'h004b,-16'h001c,-16'h0022,-16'h0005,-16'h000e,16'h0020,-16'h0021,16'h0018,-16'h002a,16'h0047,-16'h0057,16'h005c,-16'h0003,16'h0003,-16'h0020,-16'h0014,-16'h0052,-16'h0013,-16'h006f,-16'h0013,16'h0018,-16'h0010,-16'h0027,-16'h0008,-16'h0003,16'h0014,16'h005d,-16'h005f,-16'h000a,16'h0060,16'h0052,16'h0012,16'h0015,-16'h00c0,16'h0065,16'h000f,16'h0025,-16'h021f,-16'h003b,-16'h0004,-16'h0001,16'h0001,-16'h001d,16'h0008,16'h001f,16'h0010,16'h0017,16'h000e,16'h0047,16'h004c,-16'h001b,16'h0036,-16'h007e,16'h000b,-16'h0028,-16'h002d,16'h001a,16'h0029,-16'h000a,-16'h0052,16'h0027,-16'h0038,16'h004e,16'h0013,16'h0066,-16'h0011,-16'h001c,16'h005e,-16'h001a,16'h003d,-16'h0048,16'h002f,-16'h0035,16'h0045,-16'h0042,16'h0045,16'h000d,16'h0007,-16'h0017,16'h0026,-16'h0087,-16'h001d,-16'h005e,16'h000c,-16'h0004,-16'h0022,-16'h0041,16'h0002,16'h001b,16'h000c,16'h005a,-16'h0049,-16'h000d,16'h0056,16'h003f,16'h0007,16'h0011,-16'h00f4,16'h0027,-16'h0009,16'h001f,-16'h023b,-16'h0025,-16'h001c,-16'h0014,-16'h0007,-16'h0025,-16'h000d,-16'h0014,16'h001d,16'h0014,-16'h0002,16'h004e,16'h004a,-16'h001d,16'h0048,-16'h0076,-16'h0069,-16'h0028,-16'h002a,16'h0010,16'h0037,-16'h001b,-16'h001f,16'h004b,-16'h0057,16'h005c,16'h001c,16'h006c,-16'h0018,-16'h0007,16'h0066,-16'h0005,16'h002e,-16'h0086,16'h001c,-16'h001e,16'h0055,-16'h0028,16'h003e,16'h0030,16'h0010,-16'h0037,16'h0005,-16'h0049,-16'h002d,-16'h0058,-16'h0007,-16'h0013,16'h000a,-16'h0016,16'h000a,16'h0005,16'h001c,16'h0065,-16'h0076,-16'h003d,16'h0061,16'h0046,16'h0026,16'h000e,-16'h011d,-16'h0016,16'h000c,16'h0006,-16'h0220,-16'h0002,-16'h0013,16'h0004,16'h0005,-16'h0014,-16'h0003,-16'h002f,16'h001e,-16'h0002,-16'h0012,16'h004d,16'h004a,-16'h0019,16'h0032,-16'h0048,-16'h002d,16'h0016,-16'h0047,16'h000c,16'h003a,-16'h003c,16'h000e,16'h002b,-16'h0024,16'h0017,16'h0040,16'h0070,-16'h0016,16'h003f,16'h005a,16'h0008,16'h003b,-16'h00c7,16'h001e,-16'h001d,16'h0029,-16'h0038,16'h0057,16'h0023,-16'h0005,-16'h005f,-16'h0003,16'h0004,-16'h003e,-16'h0042,16'h0003,-16'h0031,16'h0011,16'h0000,16'h0024,-16'h000a,16'h0003,16'h006f,-16'h002e,-16'h0017,16'h004e,16'h0049,-16'h0002,16'h0009,-16'h012a,-16'h0025,-16'h003e,16'h0016,-16'h01fc,-16'h0019,-16'h0015,-16'h0017,16'h000b,16'h0008,-16'h000d,-16'h0004,16'h002e,-16'h000a,-16'h0032,16'h003c,16'h003a,16'h0019,16'h003b,-16'h006e,-16'h0011,16'h0023,-16'h0095,16'h0028,16'h0040,-16'h001c,16'h001a,16'h0014,-16'h001f,-16'h0041,16'h0017,16'h0069,-16'h0011,16'h0066,16'h0042,-16'h0004,16'h0031,-16'h0122,16'h0024,-16'h0040,16'h0008,-16'h0054,16'h0053,16'h0019,16'h0005,-16'h005e,-16'h0016,16'h004b,-16'h0028,-16'h0031,16'h0022,-16'h0025,-16'h0013,16'h000b,16'h000c,16'h0024,-16'h000c,16'h0063,-16'h0032,-16'h0033,16'h0050,16'h005b,16'h0000,16'h0018,-16'h0108,16'h0000,-16'h0042,16'h0035,-16'h01c2,16'h0016,16'h0003,-16'h0028,16'h0046,16'h0005,-16'h0007,-16'h0025,16'h003f,16'h0010,-16'h005a,16'h0050,16'h001d,16'h0019,16'h0001,-16'h006f,-16'h000a,16'h0041,-16'h00b3,16'h0007,16'h003e,16'h0002,16'h0057,-16'h000c,16'h0006,-16'h008b,16'h0008,16'h0061,-16'h0005,16'h0068,16'h003d,-16'h0002,16'h000e,-16'h0112,16'h0020,-16'h000f,-16'h0016,-16'h0033,16'h004d,16'h002e,-16'h0002,-16'h005a,-16'h0029,16'h004f,-16'h001c,-16'h000a,16'h002e,-16'h0051,16'h0003,-16'h000a,16'h0009,16'h002b,-16'h0002,16'h0053,-16'h0026,-16'h003b,16'h004e,16'h0051,-16'h000b,16'h001f,-16'h00c2,16'h0015,-16'h0027,16'h0023,-16'h0173,-16'h0010,16'h000a,-16'h0012,16'h0047,16'h0014,-16'h0019,-16'h0018,16'h0079,-16'h0029,-16'h0083,16'h0041,-16'h000c,16'h003c,-16'h00c2,-16'h00b0,16'h001d,16'h0040,-16'h009b,-16'h0037,16'h0023,16'h002d,16'h0064,-16'h0025,16'h0023,-16'h0050,16'h000e,16'h0035,16'h0023,16'h005a,16'h0040,16'h0000,16'h000c,-16'h00cd,16'h0021,-16'h0021,-16'h001e,-16'h0065,16'h0056,16'h002d,16'h0003,-16'h002d,-16'h0025,16'h001b,-16'h0003,16'h001c,16'h0000,-16'h0086,16'h001c,16'h0019,-16'h0001,16'h003c,-16'h006e,16'h0060,-16'h0013,-16'h0034,16'h0063,16'h0032,-16'h0010,16'h002c,-16'h0093,16'h0034,-16'h0011,16'h0032,-16'h0146,16'h0022,16'h0008,-16'h001b,16'h0018,16'h002a,-16'h003b,-16'h001b,16'h0075,-16'h002d,-16'h007b,16'h004d,-16'h001a,16'h0022,-16'h01b4,-16'h0087,16'h001e,16'h0033,-16'h0072,-16'h0058,16'h0020,16'h0069,16'h007f,-16'h0009,16'h0031,-16'h0005,16'h0000,16'h0061,16'h003a,16'h005e,16'h002c,-16'h001c,16'h0012,-16'h00ac,-16'h0003,-16'h002c,-16'h000a,-16'h004d,16'h004d,16'h0048,-16'h002b,-16'h001d,-16'h001c,16'h000b,16'h0017,16'h004e,16'h000a,-16'h00f9,16'h001a,16'h001b,-16'h001e,16'h004d,-16'h008d,16'h0055,16'h0043,-16'h001c,16'h005d,16'h0047,-16'h0010,16'h0000,-16'h0078,16'h0028,-16'h0018,16'h0012,-16'h0112,16'h001c,16'h0013,-16'h0042,-16'h000d,16'h0039,-16'h0041,-16'h001a,16'h0038,-16'h002e,-16'h00cd,16'h0053,-16'h0034,-16'h002a,-16'h01bb,-16'h00a0,16'h0026,16'h001f,-16'h0037,-16'h0059,16'h0015,16'h0083,16'h0092,-16'h0009,16'h0036,16'h003e,16'h0013,16'h006b,16'h0033,16'h0038,16'h000e,-16'h0021,16'h000a,-16'h005e,-16'h001f,-16'h0038,16'h0001,-16'h002d,16'h005b,16'h0036,-16'h0013,-16'h0048,16'h000f,-16'h002d,16'h0048,16'h0049,16'h000f,-16'h016c,16'h0025,16'h0027,-16'h0016,16'h002d,-16'h006f,16'h0057,16'h005a,-16'h001b,16'h001a,16'h0014,-16'h0016,-16'h003d,-16'h0072,16'h001a,16'h0022,16'h000a,-16'h0114,16'h0024,16'h0037,-16'h0049,-16'h0040,16'h0052,-16'h0013,-16'h0025,16'h0010,-16'h0016,-16'h00c4,16'h006c,-16'h0004,-16'h0051,-16'h0105,-16'h00b9,16'h002c,-16'h000b,-16'h0047,-16'h006c,16'h0028,16'h005d,16'h007d,16'h001d,16'h001e,16'h0031,16'h0007,16'h0054,16'h0012,16'h002c,-16'h0017,16'h0001,16'h0019,-16'h005c,16'h0010,-16'h004c,-16'h003b,16'h0041,16'h0061,16'h0034,-16'h0028,-16'h0043,-16'h000e,-16'h0068,16'h0018,16'h0053,-16'h000d,-16'h00fb,16'h0025,16'h0017,-16'h0021,-16'h0024,-16'h005b,16'h004f,16'h006b,16'h0009,16'h0045,-16'h0018,16'h0003,-16'h005f,-16'h0068,16'h0028,16'h006f,16'h0020,-16'h00ef,16'h0029,16'h0007,-16'h0022,16'h0003,16'h0040,-16'h0013,-16'h0007,16'h0014,-16'h0021,-16'h00a7,16'h008c,16'h0000,-16'h00a1,-16'h008e,-16'h0098,16'h0027,-16'h0087,-16'h002f,-16'h006a,16'h0050,16'h0022,16'h0074,16'h003b,16'h0004,16'h0044,16'h000a,16'h005a,-16'h0030,16'h003f,16'h0005,16'h0033,16'h0023,-16'h0072,16'h000b,-16'h0029,-16'h003c,16'h0068,16'h0060,16'h002b,-16'h002f,-16'h000a,-16'h0007,-16'h004c,-16'h000e,16'h0046,-16'h001d,-16'h0061,16'h002f,16'h0018,-16'h0027,-16'h0037,-16'h0058,16'h005e,16'h0021,16'h0012,16'h0011,16'h0009,16'h001a,-16'h006b,-16'h0039,-16'h001d,16'h00a8,16'h0012,-16'h00e4,16'h0021,-16'h0001,-16'h002c,16'h0036,16'h0058,16'h0007,-16'h0005,16'h000f,16'h0026,-16'h0073,16'h006a,16'h0009,-16'h008c,-16'h0024,-16'h0073,16'h002a,-16'h00e1,-16'h0004,-16'h0051,16'h0043,-16'h001b,16'h0052,16'h0021,-16'h001b,16'h002d,-16'h0016,16'h0064,-16'h0032,16'h0069,16'h0004,16'h0039,16'h0000,-16'h0060,16'h0039,-16'h0027,-16'h002a,16'h00a5,16'h0078,-16'h0003,-16'h0025,16'h0013,16'h0031,-16'h002a,-16'h0023,16'h0039,-16'h0008,-16'h003b,16'h0009,16'h0007,-16'h0025,-16'h0035,-16'h002c,16'h0053,16'h001b,-16'h001b,16'h000e,16'h0009,16'h0046,-16'h0052,-16'h0046,-16'h0033,16'h00bb,16'h002d,-16'h00ba,16'h0039,16'h0006,-16'h0032,16'h0038,16'h0052,16'h0006,16'h0010,-16'h001d,16'h0030,-16'h004b,16'h003f,-16'h0015,-16'h0043,-16'h0003,-16'h0038,16'h003d,-16'h00c0,-16'h0013,-16'h0047,-16'h000d,-16'h0024,16'h001d,16'h0029,-16'h0029,16'h003b,16'h0014,16'h0053,-16'h0043,16'h0084,-16'h0024,16'h000d,16'h0011,-16'h0036,16'h0015,-16'h0014,-16'h0013,16'h0086,16'h0059,-16'h0009,-16'h0054,16'h0025,16'h004d,-16'h0032,-16'h0034,16'h0030,-16'h0005,-16'h0021,-16'h0007,-16'h0011,16'h0003,-16'h0036,-16'h000e,16'h004f,-16'h0003,-16'h0027,16'h0011,16'h0005,16'h005a,-16'h002c,-16'h004d,-16'h002d,16'h0095,16'h0057,-16'h0089,-16'h001d,16'h0013,-16'h0032,16'h0033,16'h0072,16'h001b,16'h000f,-16'h0003,16'h0047,-16'h0030,16'h004e,-16'h0026,-16'h0003,16'h0002,-16'h0015,16'h001a,-16'h005a,16'h000b,-16'h003f,-16'h002b,16'h0022,-16'h0015,16'h0000,16'h0018,16'h003f,-16'h0015,16'h0088,-16'h003f,16'h00c2,-16'h0023,-16'h0017,-16'h0011,-16'h0028,16'h0014,-16'h001a,-16'h001a,16'h002a,16'h005f,-16'h0025,-16'h006c,-16'h000d,16'h0035,-16'h0011,-16'h0029,16'h0031,16'h000b,-16'h0002,-16'h0026,-16'h001f,16'h003f,16'h003c,16'h0021,16'h0014,16'h0001,-16'h001a,16'h003f,16'h0057,-16'h0029,16'h0041,16'h002f,16'h0023,16'h002b,-16'h0017,16'h0001,-16'h000e,-16'h0028,16'h005f,-16'h001b,16'h0009,16'h0003,-16'h0022,-16'h003a,16'h0020,16'h0041,-16'h003c,-16'h001c,-16'h0045,16'h0029,-16'h0017,16'h0000,-16'h0018,16'h0053,16'h002e,-16'h0018,-16'h0010,16'h0011,-16'h0004,16'h004b,-16'h0034,16'h0016,16'h0068,-16'h0016,16'h0000,-16'h0001,-16'h0002,16'h0003,16'h0018,16'h0005,16'h004c,16'h0042,-16'h0021,16'h0043,16'h0003,16'h000f,16'h001e,-16'h0031,-16'h0022,-16'h0029,-16'h0017,-16'h001d,16'h0005,16'h0025,-16'h0005,16'h0027,16'h0034,16'h0014,16'h001b,-16'h000d,-16'h000f,16'h0064,16'h0025,-16'h0020,16'h0034,16'h0021,16'h0027,16'h0058,-16'h002f,-16'h000e,-16'h0003,16'h0014,16'h0040,-16'h0007,16'h0000,-16'h001e,-16'h004b,-16'h0037,16'h0021,16'h0050,-16'h0022,-16'h001a,-16'h004e,16'h0027,-16'h0011,16'h001f,-16'h0005,16'h0084,16'h005a,16'h0007,16'h0000,16'h0025,-16'h001d,16'h004c,-16'h0022,16'h000b,16'h005f,-16'h0009,16'h0016,-16'h001e,-16'h000b,16'h0003,16'h002f,-16'h000b,16'h002d,16'h002b,-16'h0021,16'h004d,16'h0011,16'h000f,16'h0020,-16'h0029,-16'h0021,-16'h0040,-16'h0018,-16'h002a,-16'h0020,16'h002b,-16'h0014,16'h001f,16'h002d,16'h0006,16'h0031,-16'h000b,-16'h002e,16'h0061,16'h000e,-16'h004b,16'h004d,16'h0033,16'h0014,16'h0087,-16'h0041,-16'h0008,-16'h0020,16'h001b,16'h002d,-16'h0010,-16'h0021,-16'h001f,-16'h003f,-16'h003f,16'h0020,16'h003f,-16'h0028,-16'h0013,-16'h0046,16'h0018,-16'h0005,16'h0015,16'h0003,16'h00b2,16'h0067,16'h0036,-16'h0008,16'h001b,16'h0003,16'h0049,-16'h0034,-16'h0001,16'h0041,-16'h0018,16'h0022,-16'h0031,16'h0008,16'h0009,16'h0031,-16'h0010,16'h0032,16'h002c,-16'h004d,16'h0050,-16'h0008,16'h0010,16'h0039,-16'h0021,-16'h000c,-16'h004e,-16'h000e,-16'h0042,-16'h0016,16'h0035,-16'h000b,16'h001d,16'h0045,16'h0004,16'h003b,-16'h001a,-16'h0029,16'h006c,16'h000f,-16'h004b,16'h0040,-16'h000a,16'h0019,16'h005f,-16'h004f,-16'h002c,16'h001a,16'h0029,16'h0013,16'h000a,-16'h0030,-16'h000d,-16'h0050,-16'h0016,16'h0004,16'h0029,16'h0003,16'h0015,-16'h0069,16'h0014,16'h0000,16'h0000,-16'h0001,16'h0099,16'h005b,16'h000a,-16'h0030,16'h0042,16'h0007,16'h003d,-16'h0026,-16'h001c,16'h0050,-16'h000a,16'h000e,-16'h004f,16'h0009,-16'h000e,16'h0020,-16'h0018,16'h0013,16'h000b,-16'h004a,16'h004f,16'h0000,-16'h0004,16'h005f,-16'h0030,-16'h000d,-16'h0040,-16'h0023,-16'h003c,16'h0006,16'h000c,16'h001c,16'h0010,16'h0045,16'h001a,16'h0020,-16'h0010,-16'h0008,16'h0088,-16'h0010,-16'h0020,16'h003f,-16'h002f,-16'h0001,16'h0091,-16'h004e,-16'h0056,16'h0014,16'h0007,-16'h000b,-16'h000b,-16'h0048,-16'h0009,-16'h006a,16'h0015,-16'h0019,16'h0047,16'h0009,16'h0024,-16'h0063,16'h0019,16'h0009,-16'h0002,16'h0018,16'h009b,16'h0041,16'h001b,-16'h0034,16'h005c,-16'h0039,16'h0043,16'h0000,-16'h001b,16'h003a,-16'h0042,16'h000c,-16'h0065,16'h0025,-16'h002a,16'h0029,16'h0009,-16'h001b,16'h0008,-16'h005a,16'h0022,-16'h0018,-16'h0016,16'h001c,-16'h0038,-16'h0021,-16'h0075,-16'h0052,-16'h0017,16'h000f,16'h002e,16'h000f,16'h001c,16'h0015,16'h001c,16'h0016,-16'h0019,16'h0022,16'h0063,16'h000b,-16'h000d,16'h0019,-16'h006c,16'h000a,16'h004b,-16'h0046,-16'h0099,16'h002e,16'h0018,16'h000e,16'h0000,-16'h007b,16'h0000,-16'h004a,16'h002d,-16'h004a,16'h0011,16'h0001,16'h004f,-16'h001f,16'h003d,-16'h000b,-16'h0019,16'h0005,16'h006d,16'h002c,16'h0005,-16'h0038,16'h0062,-16'h005c,-16'h0006,16'h0019,-16'h0006,16'h0060,-16'h0032,-16'h0004,-16'h006f,16'h003d,-16'h0048,16'h001a,16'h000c,-16'h002c,-16'h0017,-16'h0037,16'h0033,-16'h0002,-16'h0030,16'h0009,-16'h001e,16'h0014,-16'h0055,-16'h008e,16'h0018,16'h0011,16'h0044,16'h000e,-16'h000a,16'h000d,16'h002f,16'h002e,-16'h0056,16'h002e,16'h006f,16'h0000,-16'h0015,16'h0032,-16'h0084,16'h0033,16'h002f,-16'h000e,-16'h00b8,16'h003d,16'h0041,16'h0017,-16'h0008,-16'h0075,-16'h000f,-16'h000e,16'h0072,-16'h002c,16'h0023,16'h001a,16'h003c,-16'h0048,16'h001b,16'h0014,-16'h006d,16'h0023,16'h004a,16'h000c,16'h000c,-16'h0034,16'h0047,-16'h008d,16'h000c,16'h0000,-16'h002f,16'h0063,16'h001a,-16'h001c,-16'h004c,16'h000b,-16'h003d,-16'h0005,-16'h0009,-16'h003f,-16'h000a,16'h0002,16'h0038,16'h0000,-16'h0010,-16'h0008,-16'h0040,-16'h0009,-16'h006d,-16'h00a6,16'h0006,16'h0038,16'h006b,16'h002e,-16'h003f,16'h0005,16'h0030,16'h0050,-16'h0084,16'h0025,16'h0064,16'h001a,16'h0004,16'h000d,-16'h00c6,16'h001f,16'h0026,16'h0018,-16'h00df,16'h0010,16'h0047,16'h0023,-16'h0023,-16'h0032,16'h001a,16'h0000,16'h0032,16'h0004,16'h002c,16'h0016,16'h0031,-16'h002a,-16'h0012,-16'h0028,-16'h0074,16'h001b,16'h003d,16'h0008,16'h0005,-16'h0013,16'h003b,-16'h006e,-16'h0007,16'h0015,-16'h0044,16'h0066,16'h003f,-16'h0029,-16'h0026,-16'h0024,-16'h0029,16'h0021,-16'h0014,-16'h003d,-16'h000f,16'h0020,16'h0039,16'h001c,-16'h0006,-16'h0026,-16'h0057,16'h002d,-16'h0066,-16'h00b4,16'h000a,16'h002c,16'h0070,16'h0002,-16'h0028,-16'h0009,16'h0017,16'h0045,-16'h00ba,16'h0043,16'h003c,16'h0039,16'h000c,16'h0001,-16'h00ac,16'h0045,16'h0019,16'h0039,-16'h0124,-16'h0003,16'h003e,16'h0012,-16'h0065,-16'h0023,16'h000d,16'h0005,16'h003d,16'h0008,16'h0030,16'h0022,-16'h0006,16'h000c,-16'h0008,-16'h0015,-16'h004e,-16'h000c,-16'h0002,-16'h0003,-16'h000c,-16'h000d,16'h001e,16'h000a,-16'h0036,16'h0008,-16'h0046,16'h0075,16'h002c,-16'h0056,-16'h001d,-16'h0037,-16'h0017,16'h0021,-16'h000a,-16'h002d,16'h000b,16'h002c,16'h004b,16'h0025,16'h0005,-16'h004e,-16'h005d,16'h002f,-16'h0074,-16'h00c6,16'h0042,16'h0049,16'h004b,-16'h0001,-16'h0013,16'h0004,-16'h0014,16'h0049,-16'h00eb,16'h0047,16'h002d,16'h0037,16'h0011,-16'h002a,-16'h00c2,16'h0062,16'h003d,16'h0035,-16'h016e,-16'h000e,16'h0042,-16'h0004,-16'h0090,-16'h003f,-16'h000d,-16'h0003,16'h0022,16'h002a,16'h0038,16'h0005,-16'h0057,16'h003b,-16'h0016,-16'h0013,-16'h0034,-16'h0021,-16'h002a,-16'h0009,-16'h0025,16'h0006,-16'h001a,16'h0015,-16'h002c,-16'h0054,-16'h000a,16'h0074,16'h000c,-16'h001e,-16'h0024,-16'h0021,-16'h0023,16'h0017,16'h0009,16'h0003,-16'h000f,16'h0044,16'h0041,16'h0033,-16'h0011,-16'h0036,-16'h0047,16'h0009,-16'h0061,-16'h009f,16'h0029,16'h0066,16'h0049,-16'h0019,-16'h0006,-16'h0008,-16'h000b,16'h005a,-16'h00d6,16'h005e,16'h0041,16'h0029,16'h0002,-16'h000b,-16'h00bb,16'h003f,16'h0023,16'h0060,-16'h018e,-16'h003e,16'h0019,16'h0007,-16'h0064,-16'h003d,16'h0024,-16'h003c,16'h001e,16'h0004,16'h0047,16'h001c,-16'h0054,16'h0028,-16'h002d,-16'h0031,16'h000d,-16'h002b,-16'h003a,-16'h0049,16'h0000,16'h0014,16'h0016,16'h0002,-16'h0032,-16'h009c,-16'h0011,16'h004f,-16'h0004,-16'h0008,-16'h0016,16'h0006,-16'h0001,16'h002c,16'h0025,16'h000e,-16'h0006,16'h0041,16'h0041,16'h0018,-16'h0002,-16'h001d,-16'h000f,16'h004a,-16'h004a,-16'h00ac,16'h0041,16'h003d,16'h0035,16'h0002,-16'h0003,-16'h0012,-16'h002c,16'h004b,-16'h00e1,16'h0048,16'h001d,16'h0033,-16'h001a,16'h0016,-16'h0092,16'h004b,-16'h0022,16'h0047,-16'h01b6,-16'h0012,16'h0015,16'h0010,-16'h0014,-16'h0051,16'h001f,-16'h002e,16'h0011,16'h001c,16'h0010,16'h000f,-16'h0032,16'h0019,-16'h0012,-16'h002f,16'h004f,-16'h0025,-16'h002b,-16'h0070,16'h0026,16'h0030,16'h0011,-16'h0032,-16'h001e,-16'h005e,-16'h0020,16'h0035,-16'h0002,16'h002d,-16'h0026,16'h000f,-16'h000a,16'h0004,16'h0009,-16'h000b,-16'h0035,16'h0021,16'h0024,16'h0000,-16'h001e,-16'h0036,-16'h000c,16'h002d,-16'h0032,-16'h00b0,16'h0024,16'h0047,16'h0009,-16'h0013,-16'h0011,16'h0002,-16'h004b,16'h002c,-16'h00c2,16'h004a,16'h0038,16'h0027,-16'h0055,16'h004e,-16'h0097,16'h0045,-16'h005d,16'h0044,-16'h01c7,-16'h0013,16'h0000,16'h0032,16'h0038,-16'h0052,16'h0025,16'h0025,16'h0016,16'h004b,16'h000d,16'h0027,-16'h001f,16'h0000,-16'h0002,-16'h0025,16'h0062,-16'h0027,-16'h002e,-16'h0054,16'h001a,-16'h0025,-16'h000c,-16'h0031,-16'h003c,-16'h005f,-16'h000d,16'h006a,16'h0001,16'h0020,-16'h0009,-16'h0014,16'h0003,-16'h0017,16'h002b,-16'h000c,-16'h0014,-16'h0010,16'h0022,16'h000e,-16'h000a,-16'h002f,16'h000d,16'h000e,-16'h0040,-16'h00e8,16'h0010,16'h004b,-16'h000f,-16'h001d,-16'h003e,16'h0021,-16'h0026,16'h003e,-16'h008c,16'h0014,16'h0028,16'h0044,-16'h0055,16'h005e,-16'h0067,16'h0048,-16'h000a,16'h0024,-16'h0187,-16'h0009,16'h0021,16'h0027,16'h0034,-16'h0080,16'h0006,16'h0030,16'h0013,16'h0028,-16'h0007,16'h0002,16'h003b,-16'h0052,-16'h0005,-16'h004b,16'h0046,-16'h002b,-16'h005c,-16'h0032,16'h0038,-16'h0027,-16'h0012,-16'h0012,-16'h0042,-16'h000b,-16'h0002,16'h0076,-16'h0016,-16'h000b,-16'h0007,-16'h0008,-16'h0003,-16'h004f,16'h0013,-16'h0011,16'h0011,-16'h0043,16'h0022,16'h0024,16'h000d,-16'h0019,16'h000a,-16'h0021,-16'h003d,-16'h0142,-16'h001b,16'h0039,-16'h003d,-16'h003d,-16'h0022,16'h0034,-16'h0013,16'h0043,-16'h0049,-16'h0003,16'h0032,16'h0054,-16'h0033,16'h004d,-16'h0085,16'h004f,16'h000c,16'h0030,-16'h0188,-16'h0013,-16'h0003,-16'h0005,16'h0052,-16'h0077,-16'h000b,16'h000e,16'h0025,16'h0019,-16'h000e,16'h0022,16'h0037,-16'h0039,16'h0023,-16'h0053,16'h0039,-16'h0005,-16'h005c,-16'h0003,16'h003e,-16'h003e,16'h0000,16'h0007,-16'h003f,16'h0025,16'h0014,16'h0091,-16'h0008,16'h0013,16'h004c,-16'h0019,16'h000c,-16'h0066,16'h0008,-16'h001f,16'h001c,-16'h0045,16'h002c,16'h000d,-16'h0004,-16'h0034,16'h0031,-16'h0057,-16'h0010,-16'h0129,-16'h0029,16'h0011,-16'h0042,-16'h001f,-16'h0022,16'h0026,16'h0018,16'h006c,-16'h0011,16'h0022,16'h0046,16'h0043,-16'h0006,16'h002f,-16'h008d,16'h0047,-16'h0007,16'h0015,-16'h017e,-16'h0026,-16'h0006,16'h0013,16'h0014,-16'h00a4,-16'h001b,-16'h000b,16'h0006,16'h0006,-16'h000d,16'h0025,16'h0063,-16'h0017,16'h0055,-16'h006a,-16'h0008,-16'h0020,-16'h0051,-16'h0004,16'h0021,-16'h0039,-16'h0016,16'h005b,-16'h0046,16'h0050,16'h001b,16'h009b,16'h0009,-16'h001d,16'h006f,-16'h001f,16'h001a,-16'h0053,-16'h000f,-16'h002f,16'h003a,-16'h004d,16'h0058,16'h0042,-16'h0009,-16'h0066,16'h0001,-16'h003f,-16'h001e,-16'h0111,-16'h0010,-16'h001b,-16'h003d,-16'h0010,-16'h000c,16'h0016,16'h000e,16'h008b,16'h0000,16'h0000,16'h0055,16'h0064,-16'h0013,16'h0014,-16'h00c0,16'h0012,16'h0022,-16'h0016,-16'h0169,16'h000f,16'h0005,-16'h0018,-16'h001e,-16'h008f,-16'h000d,-16'h000e,16'h000e,16'h0000,-16'h0011,16'h002c,16'h002e,-16'h000f,16'h004f,-16'h004c,-16'h0074,16'h0008,-16'h004e,16'h001c,16'h0057,-16'h0040,16'h0015,16'h0055,-16'h005d,16'h0057,16'h0041,16'h0090,16'h001e,16'h000b,16'h0077,-16'h001e,16'h0028,-16'h008b,16'h000b,-16'h004d,16'h0032,-16'h004c,16'h0030,16'h002e,-16'h0001,-16'h003b,16'h0021,-16'h0008,-16'h001a,-16'h00fb,-16'h000c,-16'h0033,-16'h000a,-16'h0016,16'h0023,16'h0012,16'h000d,16'h0084,-16'h0035,16'h0004,16'h002c,16'h0043,16'h0015,16'h001e,-16'h00bf,16'h0007,-16'h0010,16'h000c,-16'h0166,16'h002b,16'h0008,16'h0001,16'h0007,-16'h0089,-16'h000a,-16'h0014,16'h0018,-16'h000d,-16'h0035,16'h003b,16'h0032,-16'h003c,16'h002b,-16'h0042,-16'h0047,16'h0013,-16'h0076,16'h0009,16'h0053,-16'h003b,16'h0031,16'h006d,-16'h006b,-16'h0019,16'h002f,16'h0080,-16'h0007,16'h003c,16'h0068,-16'h0013,16'h002c,-16'h00b2,-16'h000f,-16'h002f,16'h0019,-16'h005c,16'h004d,16'h0032,-16'h0017,-16'h004e,16'h0024,16'h002c,-16'h0013,-16'h00e7,-16'h0008,-16'h0040,16'h0004,-16'h001c,16'h003a,16'h000a,16'h002e,16'h007b,-16'h0020,16'h000f,16'h003d,16'h002e,16'h002a,16'h001c,-16'h0080,-16'h001a,-16'h001e,16'h000a,-16'h0169,16'h003c,-16'h002e,-16'h0047,16'h001c,-16'h0059,-16'h0031,-16'h0043,16'h0029,16'h000f,-16'h0041,16'h004a,16'h000c,-16'h0015,16'h0034,-16'h005e,-16'h0030,16'h0033,-16'h0064,16'h0004,16'h0047,16'h0009,16'h004c,16'h0002,-16'h0044,-16'h0056,16'h002e,16'h0075,-16'h000f,16'h0055,16'h003e,16'h0000,16'h001f,-16'h00bd,-16'h000c,-16'h001f,-16'h0012,-16'h0052,16'h0053,16'h0022,16'h0011,-16'h005e,16'h0001,16'h0021,16'h000f,-16'h00c4,16'h0017,-16'h004b,16'h0007,-16'h0007,16'h004d,16'h0019,-16'h001e,16'h0061,-16'h0003,-16'h0005,16'h0049,16'h0029,16'h0005,16'h0033,-16'h0066,16'h0008,-16'h002c,16'h003b,-16'h011e,16'h0044,16'h0000,-16'h0030,16'h003d,-16'h0047,-16'h0034,-16'h0043,16'h0062,-16'h0007,-16'h004a,16'h003b,16'h0023,16'h0013,-16'h0001,-16'h0049,-16'h0022,16'h0015,-16'h006c,-16'h0010,16'h0031,16'h0042,16'h0054,-16'h0028,-16'h0009,-16'h00a9,16'h002c,16'h006a,16'h000a,16'h0071,16'h003f,-16'h000f,16'h000d,-16'h009d,16'h000d,-16'h0041,-16'h003b,-16'h004e,16'h0064,16'h0026,-16'h0024,-16'h0054,-16'h0021,16'h002f,16'h002a,-16'h00ab,16'h0002,-16'h004e,-16'h001c,16'h0001,16'h005d,16'h003f,-16'h0046,16'h0058,-16'h0013,-16'h0006,16'h0027,16'h0031,16'h000f,16'h0011,-16'h0067,-16'h001b,16'h0000,16'h0010,-16'h010d,16'h0036,16'h0007,-16'h0054,16'h0040,-16'h005c,-16'h0036,-16'h0036,16'h0094,16'h0005,-16'h007b,16'h006b,-16'h000f,16'h0017,-16'h00b8,-16'h004a,-16'h000c,16'h0025,-16'h0043,-16'h003b,16'h0034,16'h0061,16'h006d,-16'h0026,16'h001d,-16'h0075,16'h0035,16'h007f,16'h0016,16'h005a,16'h0026,-16'h000f,16'h0019,-16'h0084,16'h0017,-16'h0031,-16'h0030,-16'h0078,16'h006e,16'h0031,-16'h0034,-16'h003f,-16'h0001,16'h0027,16'h004b,-16'h0098,16'h0002,-16'h009d,16'h0018,16'h001d,16'h0034,16'h0037,-16'h0047,16'h008a,16'h0027,-16'h0001,16'h002e,16'h0035,16'h0012,16'h0015,-16'h004c,-16'h0010,16'h0024,16'h0036,-16'h0101,16'h0034,16'h0001,-16'h002d,16'h0010,-16'h003c,-16'h0064,-16'h0029,16'h008a,16'h0005,-16'h009b,16'h007d,-16'h002d,-16'h0007,-16'h0195,-16'h0040,16'h0003,16'h001d,-16'h0036,-16'h0068,16'h0022,16'h0074,16'h0069,16'h0005,16'h000b,16'h0003,16'h002a,16'h0076,16'h001a,16'h006c,-16'h0006,-16'h0020,-16'h0002,-16'h005a,16'h0009,-16'h0046,-16'h0044,-16'h004a,16'h0060,16'h0036,-16'h004d,-16'h0049,16'h0011,16'h001b,16'h0053,-16'h0067,-16'h000d,-16'h00de,16'h001e,16'h0038,16'h0027,16'h0015,-16'h0080,16'h007f,16'h005a,-16'h0003,16'h002b,16'h0038,-16'h000e,-16'h0011,-16'h006c,16'h0023,16'h0050,16'h002c,-16'h00d3,16'h0019,16'h003a,-16'h002b,-16'h002d,-16'h0031,-16'h0041,-16'h0026,16'h0075,16'h0004,-16'h008c,16'h0078,-16'h0013,-16'h0048,-16'h016f,-16'h005e,-16'h0003,16'h000b,-16'h0029,-16'h002f,16'h0033,16'h008f,16'h0053,-16'h0008,16'h0013,16'h0030,16'h0023,16'h0071,16'h001e,16'h004e,-16'h0010,-16'h000f,16'h0008,-16'h0052,16'h0000,-16'h003e,-16'h0045,-16'h0002,16'h007a,16'h0010,-16'h0066,-16'h0034,16'h000f,-16'h0038,16'h005b,-16'h0036,16'h0006,-16'h010a,16'h000a,16'h002e,16'h000e,-16'h0012,-16'h0064,16'h0045,16'h0050,16'h0009,16'h0016,16'h0000,16'h000e,-16'h0039,-16'h0043,16'h002f,16'h005b,16'h004b,-16'h00e1,16'h0022,16'h0056,-16'h0055,-16'h0047,-16'h0027,16'h000a,-16'h0037,16'h0036,16'h001f,-16'h00a5,16'h007e,16'h0016,-16'h0086,-16'h00d7,-16'h0067,16'h0018,-16'h001c,-16'h0030,-16'h003a,16'h0045,16'h0077,16'h0067,16'h0020,-16'h0002,16'h0023,16'h0024,16'h008d,-16'h002f,16'h006d,-16'h0018,16'h000a,16'h002e,-16'h005d,16'h0020,-16'h0051,-16'h003c,16'h0050,16'h00a4,-16'h0021,-16'h0077,-16'h003f,16'h001b,-16'h0065,16'h001e,-16'h0023,-16'h0001,-16'h00a0,16'h0029,16'h003c,16'h0013,-16'h0059,-16'h004c,16'h0028,16'h0068,16'h001a,16'h0021,-16'h000d,16'h0023,-16'h005e,-16'h002d,16'h0006,16'h00af,16'h0048,-16'h00d6,16'h0003,16'h0021,-16'h003a,16'h0009,-16'h0012,-16'h000b,-16'h0026,16'h0034,16'h002c,-16'h008e,16'h008a,16'h0014,-16'h0084,-16'h005e,-16'h0071,16'h002f,-16'h00a8,-16'h0015,-16'h004f,16'h0016,16'h003b,16'h006a,16'h0010,-16'h0017,16'h0046,16'h002a,16'h009f,-16'h0075,16'h0050,-16'h0020,-16'h0006,16'h000c,-16'h0054,16'h0018,-16'h0029,-16'h0041,16'h0083,16'h0066,-16'h002d,-16'h008f,-16'h002a,16'h002c,-16'h0058,-16'h004a,-16'h0030,16'h0001,-16'h0050,16'h0043,16'h0021,16'h0018,-16'h0058,-16'h0022,16'h006d,16'h0018,16'h0016,16'h002f,-16'h0005,16'h004d,-16'h004a,-16'h0035,-16'h0012,16'h00f4,16'h004b,-16'h00b3,16'h001f,-16'h000c,-16'h0017,16'h0005,16'h0005,16'h0011,-16'h0006,16'h002d,16'h0032,-16'h0078,16'h005f,16'h0005,-16'h0078,-16'h0021,-16'h004f,16'h002a,-16'h00e8,16'h0006,-16'h002d,16'h000e,16'h0037,16'h002e,16'h002d,-16'h001b,16'h0038,16'h001d,16'h00b1,-16'h007e,16'h0087,-16'h0012,-16'h0018,16'h0016,-16'h0045,16'h0039,-16'h0013,-16'h0031,16'h0065,16'h006a,-16'h0026,-16'h0052,-16'h0005,16'h006b,-16'h0043,-16'h0056,-16'h000e,-16'h0040,-16'h0007,-16'h0002,16'h0002,16'h000d,-16'h0046,-16'h000c,16'h005f,-16'h000a,-16'h0008,16'h0027,16'h0008,16'h006f,-16'h0045,-16'h0019,-16'h0023,16'h00d4,16'h0026,-16'h0095,16'h0018,-16'h0005,-16'h0024,-16'h0004,16'h000b,16'h0000,16'h0014,16'h0021,16'h0063,-16'h0063,16'h0053,-16'h0023,-16'h003f,-16'h0003,-16'h0022,16'h0012,-16'h00a1,-16'h0005,-16'h0041,-16'h0025,16'h002d,16'h002a,16'h002d,-16'h001d,16'h0012,16'h0006,16'h00c2,-16'h0065,16'h00a4,-16'h001d,-16'h003c,16'h0003,-16'h003d,16'h0021,16'h0008,-16'h000b,16'h0069,16'h0053,-16'h0021,-16'h0048,16'h0002,16'h0062,-16'h0016,-16'h0054,-16'h002a,-16'h0011,16'h000b,-16'h000f,16'h0009,16'h0018,-16'h0039,-16'h0006,16'h0050,-16'h0010,-16'h0049,16'h0012,-16'h000c,16'h0072,-16'h0034,-16'h0020,16'h0004,16'h00aa,16'h0031,-16'h0071,-16'h0007,16'h0015,-16'h0014,16'h000d,16'h006a,16'h0022,-16'h0005,16'h0008,16'h0055,-16'h0035,16'h005e,-16'h0015,-16'h000d,16'h0000,-16'h000e,16'h001c,-16'h0062,16'h0000,-16'h0014,-16'h0049,16'h002c,-16'h001a,16'h0001,16'h0012,16'h001a,-16'h000d,16'h00a2,-16'h0059,16'h00a3,-16'h001d,-16'h003b,-16'h0004,-16'h001a,16'h000d,16'h000a,-16'h0024,16'h003b,16'h0030,-16'h0038,-16'h0071,16'h000e,16'h005e,-16'h0028,-16'h004a,-16'h0012,-16'h0003,-16'h0005,-16'h002e,-16'h0019,16'h001b,16'h0015,16'h000c,16'h0000,-16'h000f,16'h0000,16'h000e,16'h0029,-16'h0003,16'h0018,16'h0014,-16'h0004,16'h001a,16'h0012,-16'h0014,-16'h0009,-16'h0010,16'h0029,-16'h000b,-16'h0011,-16'h0013,-16'h0013,-16'h0025,-16'h000a,16'h000c,-16'h0015,-16'h0006,-16'h0017,16'h0002,16'h0000,-16'h0008,-16'h0001,16'h001e,16'h0026,-16'h0004,-16'h0005,16'h0026,-16'h001e,16'h002f,-16'h0014,-16'h0001,16'h0033,16'h0012,16'h0000,-16'h0001,-16'h000c,16'h0003,16'h000c,-16'h000d,16'h0018,16'h0028,-16'h002e,16'h0028,16'h0004,16'h0025,16'h0023,16'h0000,-16'h0014,-16'h0018,-16'h0017,-16'h000d,-16'h0011,16'h0013,-16'h000a,16'h0012,16'h0020,16'h000b,16'h0008,-16'h0009,16'h0000,16'h0021,16'h0014,-16'h0012,16'h0045,16'h000e,-16'h0004,16'h0042,-16'h0006,-16'h0015,-16'h0006,-16'h0011,16'h0019,-16'h0005,16'h0002,-16'h000f,-16'h0026,-16'h0029,16'h0009,16'h003c,-16'h000e,-16'h0004,-16'h002e,16'h0002,-16'h0003,-16'h001f,-16'h0028,16'h0067,16'h0036,-16'h0008,-16'h001c,16'h0002,-16'h0001,16'h0037,-16'h0027,16'h0015,16'h0019,-16'h000b,16'h0008,-16'h001b,16'h0006,16'h0005,16'h000b,16'h0010,16'h0037,16'h0008,-16'h0035,16'h0034,-16'h0025,16'h0008,16'h0023,-16'h000d,-16'h002b,-16'h0016,-16'h0012,-16'h0019,-16'h0019,16'h0012,16'h0009,16'h001e,16'h0068,16'h0006,16'h001e,-16'h0005,-16'h0001,16'h003e,16'h0027,-16'h0029,16'h005a,-16'h0002,16'h000a,16'h0054,16'h0000,-16'h001a,-16'h0009,16'h000b,16'h002a,-16'h0027,-16'h0012,-16'h0002,-16'h0019,-16'h0007,16'h0014,16'h0030,-16'h0008,16'h0015,-16'h002e,16'h000d,16'h0001,-16'h001c,-16'h0010,16'h008a,16'h0034,16'h000c,16'h0003,16'h0034,-16'h0005,16'h0026,-16'h0001,16'h0006,16'h0042,-16'h001d,16'h0003,-16'h000d,-16'h000a,16'h0016,16'h0012,-16'h0013,16'h0015,16'h000a,-16'h001a,16'h001a,-16'h0019,-16'h0011,16'h0022,-16'h000a,-16'h0022,-16'h0036,-16'h000d,-16'h0048,-16'h0003,-16'h000b,-16'h0007,16'h0004,16'h006f,-16'h001b,16'h0026,-16'h000e,-16'h001c,16'h005a,16'h0001,-16'h0011,16'h006b,-16'h0024,16'h000f,16'h0049,-16'h0026,-16'h0031,16'h000b,16'h0010,16'h000e,-16'h0013,-16'h0019,-16'h0022,-16'h004f,-16'h0002,-16'h0009,16'h005a,-16'h0013,16'h0006,-16'h002e,-16'h0018,-16'h0004,-16'h001a,16'h0005,16'h008b,16'h0041,-16'h0006,-16'h001c,16'h0041,-16'h0016,16'h0051,16'h0008,-16'h000a,16'h002c,-16'h000b,16'h000c,-16'h0019,16'h0009,16'h0000,16'h0012,-16'h001f,16'h000f,16'h0014,-16'h0021,16'h0036,-16'h0004,-16'h002b,16'h0015,-16'h002e,-16'h0011,-16'h0033,-16'h0009,-16'h0041,-16'h0011,16'h000e,16'h0012,-16'h0004,16'h0048,16'h000e,16'h001c,-16'h0015,16'h0021,16'h005b,16'h0002,-16'h003b,16'h0059,-16'h004d,16'h0003,16'h005c,-16'h0021,-16'h002d,16'h0015,-16'h0006,16'h0011,-16'h0038,-16'h0018,-16'h0014,-16'h0039,16'h000b,-16'h0016,16'h004a,-16'h0017,16'h002a,-16'h0020,-16'h0002,16'h0010,-16'h0029,16'h001d,16'h0097,16'h0020,16'h0017,-16'h0039,16'h005f,-16'h0003,16'h004c,-16'h0003,16'h0005,16'h0012,-16'h001c,16'h0027,-16'h004f,16'h001a,-16'h001d,16'h001e,16'h0003,-16'h0019,-16'h0005,-16'h0037,16'h0023,-16'h0015,-16'h0021,16'h0002,-16'h0034,-16'h0026,-16'h005d,-16'h0039,-16'h002f,16'h0012,16'h0021,16'h001a,-16'h0005,16'h0069,16'h0001,16'h0023,-16'h002b,16'h002e,16'h0050,-16'h000b,-16'h000e,16'h0047,-16'h0050,-16'h0003,16'h0052,-16'h0015,-16'h005f,16'h0049,16'h0017,16'h0028,-16'h0041,-16'h004b,-16'h0011,-16'h0018,16'h0017,-16'h0036,16'h003d,-16'h000b,16'h0031,-16'h003b,16'h0025,16'h0002,-16'h005d,16'h0017,16'h009d,16'h001a,-16'h0008,-16'h002d,16'h0032,-16'h001c,16'h002e,-16'h0003,-16'h0014,16'h001c,-16'h001a,16'h0014,-16'h0049,16'h0017,-16'h002d,16'h002b,16'h0000,-16'h0025,-16'h0002,-16'h0021,16'h0018,-16'h0002,-16'h000f,-16'h000a,-16'h005f,-16'h0009,-16'h004f,-16'h004a,-16'h0006,16'h001b,16'h0038,16'h000d,-16'h0016,16'h0032,16'h0036,16'h0015,-16'h002c,16'h0045,16'h003e,-16'h0023,16'h0001,16'h004e,-16'h0079,16'h0010,16'h005b,-16'h0023,-16'h008b,16'h003b,16'h0027,16'h0021,-16'h004a,-16'h0039,16'h000d,16'h0006,16'h002b,-16'h0026,16'h004d,-16'h0001,16'h0054,-16'h0027,-16'h0006,16'h001e,-16'h008a,-16'h0005,16'h005b,16'h000a,16'h0004,-16'h000c,16'h001c,-16'h0022,16'h0031,16'h000b,-16'h0012,16'h0045,16'h0021,16'h000a,-16'h0056,16'h0013,-16'h002f,16'h0024,-16'h0022,-16'h004b,16'h0014,-16'h0013,16'h000c,16'h0010,-16'h002d,-16'h000b,-16'h0069,16'h0022,-16'h0072,-16'h0079,16'h0009,16'h003a,16'h006f,16'h0010,-16'h0014,16'h0016,16'h003b,16'h000e,-16'h0053,16'h0033,16'h0040,-16'h0012,16'h000a,16'h0013,-16'h0089,16'h000d,16'h0048,16'h0017,-16'h00aa,16'h001f,16'h002e,16'h003f,-16'h0042,-16'h002d,16'h000b,16'h000a,16'h002b,-16'h0010,16'h004a,-16'h0004,16'h0037,-16'h0030,16'h0009,-16'h0002,-16'h005d,-16'h0008,-16'h000a,16'h0005,16'h0003,-16'h001a,16'h0016,-16'h0011,16'h0006,-16'h000a,-16'h0030,16'h002f,16'h0044,-16'h0031,-16'h0016,16'h0006,-16'h0021,16'h0030,-16'h0020,-16'h004f,-16'h0008,-16'h000d,16'h0024,16'h0019,16'h0000,-16'h0021,-16'h0073,16'h0028,-16'h0078,-16'h006f,-16'h0009,16'h002b,16'h005f,16'h001a,-16'h0015,16'h0027,16'h001d,16'h000e,-16'h0074,16'h003f,16'h0032,-16'h000b,16'h0016,16'h0005,-16'h0079,16'h0046,16'h004c,16'h0036,-16'h009c,-16'h0012,16'h0031,16'h0036,-16'h0099,16'h0007,16'h001d,16'h0025,16'h002c,16'h0009,16'h0044,-16'h000c,-16'h002c,16'h0000,-16'h002a,-16'h0007,-16'h0055,-16'h002d,-16'h0024,16'h000c,-16'h0008,-16'h0012,-16'h000e,16'h001d,-16'h0030,-16'h0024,-16'h0030,16'h002f,16'h0022,-16'h0034,16'h0000,-16'h0007,-16'h0032,16'h003a,16'h0019,-16'h0024,-16'h0021,16'h0008,16'h0027,16'h001c,16'h0006,-16'h0028,-16'h0061,16'h0019,-16'h0065,-16'h006c,16'h002d,16'h0035,16'h003e,16'h0017,-16'h0004,16'h002e,-16'h0012,16'h001e,-16'h005a,16'h0055,16'h0038,-16'h0002,16'h001d,-16'h000a,-16'h0092,16'h0054,16'h002f,16'h0041,-16'h00c5,-16'h0032,16'h0014,16'h0014,-16'h00a5,-16'h0009,16'h0039,-16'h0003,16'h0022,16'h0032,16'h0048,16'h0000,-16'h0066,16'h002d,-16'h0014,-16'h0033,-16'h0011,-16'h0028,-16'h0021,-16'h0018,-16'h0022,-16'h0026,16'h0008,16'h000d,-16'h0022,-16'h0081,-16'h0032,16'h0053,-16'h0005,-16'h0030,16'h0025,-16'h003f,-16'h001d,16'h0017,16'h0014,-16'h0021,-16'h0020,16'h0015,16'h0032,16'h0014,-16'h0016,-16'h004d,-16'h005b,16'h002b,-16'h0052,-16'h0066,16'h0038,16'h0051,16'h0029,16'h000d,-16'h0031,-16'h0015,-16'h002e,16'h001a,-16'h0077,16'h0059,16'h0036,16'h000b,16'h0022,16'h0003,-16'h007b,16'h005b,16'h002c,16'h0062,-16'h00cd,-16'h0037,16'h0004,16'h0025,-16'h0045,-16'h000e,16'h0035,-16'h0022,16'h001c,16'h0021,16'h0035,16'h0003,-16'h006d,16'h0015,-16'h0008,-16'h001f,16'h0052,-16'h002d,-16'h0053,-16'h005b,16'h0019,16'h0003,16'h0009,-16'h0017,-16'h0021,-16'h0061,-16'h001a,16'h0041,-16'h002c,-16'h0004,16'h0016,-16'h000a,-16'h0012,16'h0009,16'h0012,-16'h0026,-16'h0008,16'h0024,16'h0026,16'h0034,-16'h0019,-16'h003f,-16'h003c,16'h0025,-16'h0062,-16'h0064,16'h0041,16'h0020,16'h000d,16'h0034,-16'h0033,-16'h000d,-16'h005a,16'h001f,-16'h0060,16'h0035,16'h000f,16'h0000,-16'h0023,16'h001b,-16'h0085,16'h003a,-16'h002c,16'h005f,-16'h00d1,-16'h0028,-16'h0016,16'h0012,16'h001a,-16'h0017,16'h002d,-16'h0031,16'h002f,16'h0025,16'h0020,16'h000b,-16'h005f,-16'h000c,-16'h001d,-16'h0027,16'h006e,-16'h0010,-16'h0040,-16'h006c,16'h0021,16'h000e,16'h0015,-16'h0043,-16'h002c,-16'h0047,-16'h002f,16'h0048,-16'h0015,-16'h0018,16'h004b,-16'h000f,-16'h0013,-16'h001e,16'h000d,-16'h001c,-16'h0035,16'h0034,16'h0046,16'h0007,-16'h002c,-16'h0035,-16'h0020,-16'h000f,-16'h004c,-16'h006a,16'h0000,16'h0010,-16'h0028,-16'h0003,-16'h0023,16'h000b,-16'h0059,16'h0022,-16'h004b,16'h002c,16'h0008,16'h0004,-16'h003c,16'h0041,-16'h007f,16'h0021,-16'h0029,16'h003a,-16'h00cc,16'h0008,16'h0015,16'h0022,16'h0040,-16'h0008,16'h002e,16'h0003,16'h002f,16'h004c,-16'h0008,16'h0007,-16'h0011,16'h0000,-16'h000e,-16'h0025,16'h0076,-16'h001d,-16'h0062,-16'h004d,16'h002f,-16'h0036,-16'h0007,-16'h0019,-16'h0047,16'h0007,-16'h0016,16'h0038,-16'h000c,16'h0026,16'h0045,-16'h0018,16'h0002,-16'h0049,16'h0009,16'h0010,-16'h003a,-16'h0013,16'h001f,16'h0013,-16'h0011,-16'h002a,16'h0011,-16'h0016,-16'h001e,-16'h0096,-16'h0011,16'h0024,-16'h0036,-16'h001e,-16'h001d,16'h0039,-16'h0039,16'h002f,-16'h0047,16'h0001,16'h0024,16'h0022,-16'h0041,16'h004e,-16'h005a,16'h0033,-16'h003b,16'h0010,-16'h00ea,16'h0014,16'h0019,16'h0020,16'h004f,-16'h0020,16'h0005,16'h000b,16'h002b,16'h0052,-16'h003a,16'h0020,16'h002c,-16'h002a,-16'h0002,-16'h0028,16'h005d,-16'h0009,-16'h0099,-16'h0043,16'h0034,-16'h0055,16'h0019,-16'h0007,-16'h0054,16'h0018,-16'h001f,16'h0074,-16'h000a,16'h0021,16'h0055,-16'h0028,-16'h0018,-16'h0074,16'h001f,16'h0002,-16'h000d,-16'h0026,16'h0039,16'h0014,-16'h001b,-16'h0019,16'h003e,-16'h0038,-16'h0022,-16'h00c1,-16'h0004,16'h001f,-16'h0032,-16'h0017,-16'h0011,16'h003b,-16'h000b,16'h002d,-16'h0011,16'h0019,16'h001f,16'h0044,-16'h0044,16'h003b,-16'h0071,16'h0023,-16'h0005,16'h0015,-16'h00d2,-16'h0009,-16'h000b,16'h0019,16'h0046,-16'h0047,16'h0011,16'h0014,16'h0051,16'h002d,-16'h0044,16'h0015,16'h0049,-16'h0035,16'h0024,-16'h0022,16'h0040,16'h001f,-16'h007f,-16'h001a,16'h003d,-16'h0057,-16'h0006,16'h0003,-16'h005b,16'h0065,-16'h0003,16'h0071,-16'h0009,-16'h0007,16'h0069,-16'h000d,-16'h0003,-16'h0075,16'h0009,16'h0000,16'h0000,-16'h0079,16'h004c,16'h001f,-16'h0012,-16'h004f,16'h0037,-16'h0059,-16'h0009,-16'h00f6,-16'h000b,-16'h000e,-16'h0049,-16'h002b,-16'h0017,16'h0045,-16'h001f,16'h0052,-16'h0001,16'h003d,-16'h0015,16'h0055,-16'h0005,16'h0017,-16'h0063,16'h001d,16'h0008,-16'h000a,-16'h00c0,16'h0016,16'h0009,-16'h002d,16'h0026,-16'h0052,-16'h0026,-16'h000e,16'h0039,16'h0009,-16'h0056,16'h0018,16'h003f,-16'h0032,16'h0012,-16'h003e,16'h0011,16'h0015,-16'h0089,16'h0016,16'h0051,-16'h0054,16'h000b,16'h0048,-16'h0055,16'h0052,16'h000a,16'h007e,16'h0004,-16'h0013,16'h0060,-16'h0009,16'h003a,-16'h007f,16'h000c,-16'h0016,16'h000b,-16'h0084,16'h0061,16'h0024,-16'h0020,-16'h0063,16'h0033,-16'h0026,-16'h0007,-16'h012b,16'h0009,-16'h0055,-16'h004d,-16'h002c,-16'h0008,16'h002d,16'h0015,16'h0074,16'h0016,16'h002e,16'h000f,16'h0047,-16'h001a,16'h0020,-16'h0053,16'h001f,16'h0011,-16'h0030,-16'h00b5,16'h0020,16'h0005,-16'h0021,16'h000b,-16'h0077,-16'h0015,-16'h0016,16'h000e,16'h0006,-16'h0032,16'h0000,16'h001a,-16'h0038,16'h0033,-16'h0027,-16'h0077,16'h0007,-16'h0044,16'h0032,16'h0048,-16'h0056,16'h002a,16'h0077,-16'h003c,16'h0015,16'h0028,16'h0099,16'h0013,-16'h0005,16'h0098,-16'h002d,16'h003b,-16'h0081,16'h0005,16'h0008,16'h001d,-16'h0080,16'h005b,16'h003a,-16'h0015,-16'h005b,16'h0033,-16'h0008,-16'h0001,-16'h0153,16'h000d,-16'h0057,-16'h001f,-16'h0033,-16'h0009,16'h0015,-16'h0003,16'h007a,16'h0010,16'h002a,16'h001b,16'h003a,-16'h0010,16'h001a,-16'h0042,16'h000d,16'h001e,-16'h001d,-16'h00ca,16'h0022,-16'h0001,-16'h002a,16'h0012,-16'h008c,-16'h003b,-16'h0022,16'h000e,16'h0005,-16'h0063,16'h0018,-16'h0001,-16'h005d,16'h0006,-16'h0028,-16'h003a,16'h0031,-16'h0024,16'h0035,16'h0067,-16'h0026,16'h0050,16'h0047,-16'h006f,-16'h0011,16'h0034,16'h006a,16'h001f,16'h001c,16'h0038,16'h0006,16'h001c,-16'h0077,16'h0003,-16'h0017,-16'h0022,-16'h0063,16'h0066,16'h0034,-16'h000e,-16'h0085,16'h0025,16'h001c,16'h001d,-16'h015c,-16'h0017,-16'h002c,16'h001d,-16'h000f,16'h0006,16'h002d,-16'h0023,16'h007e,16'h001a,16'h0031,16'h004d,16'h005c,-16'h0016,16'h0016,-16'h0033,16'h000b,-16'h000a,-16'h0015,-16'h00a8,16'h004a,-16'h000b,-16'h0073,16'h004d,-16'h0097,-16'h0052,-16'h0013,16'h0011,-16'h0027,-16'h0054,16'h0033,16'h0011,-16'h0029,16'h0021,-16'h002d,-16'h001e,16'h0013,-16'h0030,-16'h0001,16'h003b,16'h000a,16'h0046,16'h0000,-16'h0049,-16'h006e,16'h001b,16'h0070,16'h000c,16'h0037,16'h004f,16'h0008,16'h001c,-16'h0080,16'h0010,-16'h0005,-16'h0031,-16'h005f,16'h005e,16'h0036,-16'h0014,-16'h0061,16'h0021,16'h0052,16'h001e,-16'h016f,-16'h0001,-16'h0050,16'h001c,-16'h0012,-16'h0006,16'h0033,-16'h0055,16'h009c,16'h0013,16'h001e,16'h0026,16'h003e,-16'h003a,16'h0017,-16'h0028,-16'h001c,16'h0005,16'h000b,-16'h00c3,16'h0068,-16'h0018,-16'h0091,16'h004f,-16'h009a,-16'h0058,-16'h003f,16'h004c,-16'h0013,-16'h0035,16'h0037,-16'h001c,-16'h001d,-16'h0025,-16'h001b,-16'h002f,16'h0020,-16'h000b,-16'h000c,16'h0030,16'h003b,16'h0064,-16'h003c,-16'h000e,-16'h0094,16'h0030,16'h006e,16'h0020,16'h005b,16'h003d,16'h0005,16'h001c,-16'h0074,16'h000f,-16'h0033,-16'h0012,-16'h004c,16'h0082,16'h0025,-16'h0045,-16'h005a,-16'h001f,16'h004d,16'h0043,-16'h0135,-16'h0024,-16'h005b,16'h0005,-16'h0004,16'h0010,16'h0027,-16'h0079,16'h0074,16'h0016,-16'h0015,16'h003a,16'h0009,-16'h0023,16'h0018,-16'h0034,-16'h0021,16'h000a,16'h0028,-16'h00de,16'h004a,-16'h0001,-16'h0046,16'h0056,-16'h00a4,-16'h0052,-16'h0067,16'h00a6,-16'h0013,-16'h0066,16'h0044,-16'h0025,16'h0000,-16'h00bb,-16'h0023,-16'h0011,16'h0027,-16'h001b,-16'h0027,16'h0037,16'h0076,16'h0061,-16'h001c,-16'h0003,-16'h005e,16'h004a,16'h008c,16'h0012,16'h0068,16'h000c,16'h0000,16'h001a,-16'h0075,16'h0035,-16'h002c,-16'h0050,-16'h0077,16'h005a,16'h0021,-16'h008c,-16'h0066,16'h0014,16'h0030,16'h0049,-16'h0101,-16'h0022,-16'h00a5,-16'h000b,16'h000f,16'h003a,16'h0005,-16'h0069,16'h0090,16'h002f,16'h0003,16'h0049,16'h001e,-16'h0021,-16'h000c,-16'h003a,-16'h0021,16'h0058,16'h0044,-16'h00cd,16'h000d,16'h0000,-16'h0056,16'h0000,-16'h00a9,-16'h002e,-16'h0043,16'h0091,16'h000d,-16'h007c,16'h003f,-16'h000f,-16'h0008,-16'h015c,-16'h0017,16'h0006,16'h0000,-16'h0020,-16'h002d,16'h003f,16'h007d,16'h0064,-16'h000f,-16'h0011,-16'h000e,16'h0041,16'h0093,-16'h0020,16'h0065,16'h0024,-16'h0026,16'h0009,-16'h0061,16'h0017,-16'h0046,-16'h0037,-16'h004e,16'h006f,16'h000f,-16'h0070,-16'h005c,16'h002e,16'h0005,16'h003d,-16'h00e6,-16'h0020,-16'h00ca,16'h0022,16'h0035,16'h0048,-16'h000e,-16'h004c,16'h0062,16'h0038,-16'h0005,16'h0045,16'h0011,-16'h0008,-16'h002a,-16'h003c,16'h000a,16'h0063,16'h005c,-16'h00ae,16'h0018,16'h001a,-16'h0057,-16'h0028,-16'h00a2,-16'h0014,-16'h0040,16'h0072,16'h0027,-16'h0093,16'h005f,-16'h001c,-16'h0041,-16'h0111,-16'h0007,-16'h0001,16'h0017,-16'h001d,-16'h0045,16'h0045,16'h007c,16'h007c,16'h000e,16'h0018,16'h0022,16'h0047,16'h00be,-16'h0017,16'h006d,16'h0013,-16'h004a,16'h0019,-16'h0055,16'h0024,-16'h002d,-16'h002c,16'h000f,16'h006f,-16'h0011,-16'h008b,-16'h004e,16'h003d,-16'h001e,16'h0036,-16'h00af,-16'h0020,-16'h00cd,16'h0035,16'h002a,16'h003f,-16'h0031,-16'h002d,16'h000c,16'h004e,16'h0011,16'h000d,-16'h0024,16'h0031,-16'h0056,-16'h0017,16'h0021,16'h007f,16'h0036,-16'h00c2,-16'h0001,16'h0017,-16'h006d,-16'h003c,-16'h005d,16'h000a,-16'h004e,16'h004f,16'h003f,-16'h0089,16'h0064,-16'h0024,-16'h0076,-16'h0092,-16'h002e,16'h001d,-16'h0028,-16'h000c,-16'h003b,16'h0055,16'h0068,16'h0077,16'h0003,16'h002a,16'h001b,16'h005d,16'h00ac,-16'h0050,16'h0055,-16'h0018,-16'h0027,16'h001d,-16'h003d,16'h0029,-16'h000f,-16'h0032,16'h0052,16'h0058,-16'h001d,-16'h0096,-16'h0043,16'h0032,-16'h003e,-16'h0025,-16'h00a0,16'h0005,-16'h0085,16'h0041,16'h002e,16'h0023,-16'h0062,-16'h0003,16'h0032,16'h002b,16'h0025,16'h0026,-16'h000d,16'h0031,-16'h004b,-16'h0005,16'h001a,16'h00cb,16'h0059,-16'h00ad,16'h000f,16'h0020,-16'h0034,-16'h000a,-16'h0052,16'h0003,-16'h0027,16'h004e,16'h002d,-16'h007c,16'h0052,-16'h000f,-16'h0072,-16'h0046,-16'h0022,16'h0021,-16'h007c,16'h0009,-16'h0062,16'h0049,16'h006f,16'h008b,16'h0003,16'h0020,16'h0054,16'h0043,16'h00d5,-16'h0088,16'h004c,16'h0000,-16'h000f,16'h001c,-16'h0036,16'h0010,-16'h0006,-16'h0038,16'h0054,16'h0056,-16'h001e,-16'h006f,-16'h0003,16'h0054,-16'h0049,-16'h004c,-16'h0093,16'h0006,-16'h0044,16'h003e,16'h0043,16'h0034,-16'h006e,-16'h0006,16'h003a,16'h0008,16'h0003,16'h003b,-16'h002e,16'h0060,-16'h0037,-16'h0017,-16'h0020,16'h00c6,16'h0027,-16'h008f,16'h004f,-16'h000f,-16'h0028,16'h000c,-16'h003e,16'h0016,-16'h0009,16'h0040,16'h0059,-16'h0059,16'h0041,-16'h0019,-16'h004d,-16'h000d,-16'h000c,16'h000f,-16'h009f,-16'h0012,-16'h0032,-16'h0007,16'h001e,16'h0069,16'h0035,-16'h0014,16'h0039,16'h002a,16'h00c9,-16'h0078,16'h006f,-16'h0019,-16'h0041,16'h0017,-16'h0022,16'h000e,16'h0022,-16'h002d,16'h008f,16'h0036,-16'h0031,-16'h0053,-16'h0004,16'h0060,-16'h003b,-16'h0041,-16'h008f,-16'h001a,-16'h0014,16'h0022,16'h0048,16'h0039,-16'h0060,16'h000a,16'h0023,16'h0002,-16'h000b,16'h0013,16'h0008,16'h007d,-16'h0022,-16'h0010,-16'h0020,16'h00c4,16'h0043,-16'h0092,16'h000c,16'h0015,-16'h001e,-16'h000e,-16'h000a,16'h002e,16'h000d,16'h0033,16'h0046,-16'h0032,16'h0040,-16'h0021,-16'h001d,16'h0000,-16'h000a,16'h0012,-16'h0075,-16'h0002,-16'h001d,-16'h001f,16'h003d,16'h0000,16'h0019,16'h0004,16'h0009,-16'h000e,16'h00b5,-16'h0076,16'h0072,-16'h0021,-16'h0042,-16'h001c,-16'h002a,16'h0014,-16'h0009,-16'h000a,16'h005f,16'h001f,-16'h003a,-16'h0033,16'h001b,16'h007c,-16'h0020,-16'h004b,-16'h0052,-16'h0013,16'h000b,-16'h001e,16'h0005,16'h0014,-16'h0024,16'h0018,16'h0027,16'h0016,-16'h001c,16'h000e,16'h0008,16'h0078,-16'h0002,16'h000a,16'h0007,16'h0085,16'h0038,-16'h0071,-16'h0031,-16'h0003,-16'h0004,-16'h0008,16'h001e,16'h0020,16'h0012,16'h000f,16'h002b,-16'h0020,16'h0029,-16'h003d,16'h0001,-16'h0005,16'h000e,-16'h0018,-16'h0036,-16'h0006,-16'h000f,-16'h004e,16'h0016,-16'h000c,-16'h0001,16'h0014,16'h0001,-16'h0022,16'h0095,-16'h0046,16'h0096,-16'h0013,-16'h003a,-16'h003a,-16'h0011,16'h001d,-16'h0020,-16'h0018,16'h003a,16'h0030,-16'h0020,-16'h0046,16'h0005,16'h0046,-16'h0031,-16'h0040,-16'h003a,16'h0006,16'h001c,-16'h0022,-16'h001c,16'h0001,16'h0008,16'h0000,-16'h000f,16'h0004,-16'h0003,-16'h0004,16'h0003,16'h0000,16'h0004,-16'h000a,-16'h000a,16'h0006,16'h0000,-16'h0008,16'h0009,-16'h0001,16'h001d,-16'h0007,16'h000d,-16'h0008,-16'h001a,-16'h000b,16'h0000,-16'h0005,16'h0003,16'h000a,-16'h000d,16'h0007,-16'h0004,-16'h0006,-16'h0011,16'h000f,16'h0000,-16'h0006,-16'h0003,16'h0009,16'h000d,16'h0015,-16'h0016,16'h000c,16'h000c,16'h000c,-16'h0001,-16'h0009,-16'h000d,16'h000e,16'h0014,16'h000a,16'h001e,16'h0005,16'h0003,16'h0009,16'h0002,16'h0017,16'h0003,-16'h0007,-16'h000d,-16'h0019,16'h0005,-16'h0003,16'h0016,16'h0011,-16'h0018,-16'h0001,16'h0016,-16'h0007,16'h000a,-16'h0013,-16'h000c,-16'h0008,16'h0015,16'h000b,16'h0017,-16'h0007,16'h0008,16'h0025,-16'h0001,-16'h0006,16'h0001,-16'h0013,-16'h0002,-16'h0009,16'h000c,-16'h000f,-16'h0003,-16'h000f,16'h0002,16'h000c,-16'h0014,16'h0012,-16'h001c,-16'h0013,-16'h0004,-16'h000d,16'h0003,16'h0044,16'h0021,16'h000d,-16'h000e,16'h0013,-16'h0004,16'h0021,16'h0000,16'h000f,16'h000e,16'h0012,-16'h0003,16'h0001,16'h0003,16'h0005,-16'h000d,16'h000d,16'h0002,16'h0016,-16'h0016,16'h0000,-16'h0021,16'h0002,16'h000f,16'h0001,-16'h001e,-16'h0005,16'h0007,16'h0003,16'h000b,-16'h0012,16'h0000,16'h001e,16'h0026,-16'h000e,16'h0004,-16'h000a,-16'h0001,-16'h0003,16'h0001,-16'h0008,16'h0024,-16'h0008,16'h0004,16'h0021,16'h0019,16'h0010,-16'h0018,16'h001a,-16'h0004,-16'h0001,16'h0000,16'h0004,-16'h0001,-16'h000f,-16'h0007,16'h000b,-16'h0005,16'h0010,-16'h0024,16'h0009,16'h0000,-16'h000c,-16'h001e,16'h0063,16'h0027,16'h0013,16'h0002,16'h0012,-16'h000c,16'h002c,-16'h0016,16'h000f,16'h0009,16'h0002,16'h001a,-16'h001b,16'h0020,16'h0001,16'h0007,-16'h0001,16'h0028,-16'h000a,-16'h0014,16'h0000,-16'h0006,-16'h0014,16'h0029,-16'h0008,-16'h0013,-16'h0025,-16'h0004,-16'h0016,16'h0014,-16'h0003,-16'h0010,-16'h0012,16'h0038,-16'h000a,16'h0003,-16'h0018,-16'h0006,16'h001a,16'h0000,-16'h001c,16'h003d,-16'h0029,-16'h0002,16'h0021,16'h000f,-16'h000b,-16'h000c,-16'h0003,16'h001d,-16'h000e,-16'h0015,16'h0000,-16'h0013,-16'h0006,-16'h000e,16'h0034,16'h0003,16'h0027,-16'h002e,-16'h0011,-16'h0007,-16'h002a,16'h000a,16'h0068,16'h0024,-16'h0002,-16'h0017,16'h0007,16'h0000,16'h002c,16'h0009,16'h0002,16'h0010,-16'h0018,16'h000d,-16'h0029,16'h002c,16'h001a,16'h001c,-16'h000d,16'h001e,16'h0013,-16'h0032,16'h0002,-16'h0013,-16'h0025,16'h0021,-16'h000a,-16'h0010,-16'h0019,-16'h0014,-16'h0039,-16'h000d,16'h0001,-16'h000f,-16'h0006,16'h0041,-16'h0007,16'h0005,16'h0008,16'h000f,16'h002b,-16'h0025,-16'h001a,16'h0042,-16'h002a,-16'h0033,16'h002b,-16'h0007,-16'h001e,16'h002a,16'h0003,16'h0030,-16'h0011,-16'h0016,-16'h001c,-16'h0014,16'h0005,-16'h0016,16'h0065,16'h0008,16'h0042,-16'h001a,-16'h0005,-16'h0003,-16'h0032,16'h001c,16'h0066,16'h0046,16'h0017,16'h0000,16'h0015,16'h0001,16'h0032,16'h0013,16'h0016,16'h0003,-16'h0014,16'h0028,-16'h0028,16'h002c,16'h000a,16'h0019,-16'h0001,16'h001f,-16'h0020,-16'h003a,16'h001d,16'h000a,-16'h001d,-16'h000c,-16'h003d,-16'h0004,-16'h0047,-16'h0026,-16'h0036,16'h001c,16'h0006,-16'h0024,-16'h0031,16'h005a,16'h0001,16'h0008,-16'h0029,16'h0004,16'h000f,-16'h002f,-16'h003c,16'h0045,-16'h004d,-16'h000e,16'h0050,16'h0015,-16'h0036,16'h0040,16'h0002,16'h001f,-16'h0033,-16'h0027,-16'h0014,-16'h0030,-16'h0012,-16'h0003,16'h0047,-16'h0007,16'h004b,-16'h0025,16'h0007,-16'h0009,-16'h0063,16'h000b,16'h0052,16'h0044,-16'h0001,16'h0019,16'h0019,16'h0023,16'h0059,16'h0000,-16'h000e,16'h0015,-16'h0023,16'h0007,-16'h0043,16'h0040,-16'h0026,16'h002e,-16'h001c,16'h0015,-16'h0008,-16'h0024,16'h000e,-16'h0001,-16'h004c,-16'h0004,-16'h0050,16'h0008,-16'h0044,-16'h001e,-16'h001a,16'h0046,-16'h0005,-16'h0016,-16'h000f,16'h0060,16'h0007,16'h0006,-16'h0012,16'h0021,16'h0014,-16'h003a,-16'h0028,16'h0018,-16'h005b,-16'h000d,16'h0033,16'h0016,-16'h0052,16'h0058,16'h0000,16'h0018,-16'h0040,-16'h0014,-16'h001c,-16'h0017,-16'h0033,-16'h001a,16'h0052,-16'h0006,16'h005a,-16'h0008,-16'h0023,16'h0014,-16'h0071,-16'h0007,16'h0045,16'h0044,-16'h0018,16'h0009,-16'h0006,16'h0037,16'h0042,16'h000d,-16'h001f,16'h0030,16'h0017,16'h0010,-16'h0042,16'h0009,-16'h004a,16'h004e,-16'h0020,-16'h0002,-16'h0035,-16'h003b,16'h0009,-16'h0006,-16'h003e,-16'h0023,-16'h0073,16'h003d,-16'h0035,-16'h002c,-16'h0041,16'h006e,16'h0004,-16'h002e,-16'h0030,16'h0057,16'h001a,-16'h0003,-16'h001e,16'h0027,16'h002f,-16'h001f,-16'h0024,16'h0016,-16'h004d,16'h0014,16'h004f,16'h0040,-16'h0071,16'h003a,-16'h0003,16'h0035,-16'h0064,-16'h001b,-16'h000d,-16'h0034,-16'h001f,16'h0000,16'h0055,-16'h0019,16'h004b,-16'h0010,-16'h003d,-16'h0008,-16'h0053,-16'h0003,16'h000d,16'h0055,-16'h0006,16'h0006,-16'h0012,16'h0042,16'h0010,16'h0011,-16'h0020,16'h0046,16'h0028,16'h0005,-16'h0017,-16'h0005,-16'h0034,16'h0053,16'h0007,16'h0000,-16'h0039,-16'h0062,16'h001f,-16'h0008,-16'h0034,-16'h0018,-16'h008c,16'h0053,-16'h005e,-16'h0035,-16'h0037,16'h007a,16'h0021,-16'h0021,16'h0002,16'h004a,16'h0009,-16'h0029,-16'h0020,16'h0016,16'h0025,-16'h0022,-16'h0004,16'h0007,-16'h0055,16'h0042,16'h0036,16'h0058,-16'h0068,16'h0002,-16'h0011,16'h0025,-16'h0095,16'h0022,16'h0004,-16'h001f,-16'h0017,16'h000f,16'h0084,-16'h001b,-16'h0013,-16'h0003,-16'h003d,16'h0010,-16'h003b,-16'h0008,-16'h000a,16'h0021,-16'h0003,-16'h0015,16'h000e,16'h004c,-16'h0004,-16'h0031,-16'h0023,16'h002e,16'h002b,-16'h001d,16'h0011,-16'h001a,-16'h0034,16'h006e,-16'h0009,-16'h0017,-16'h0032,-16'h0058,16'h0044,16'h0008,-16'h0043,-16'h002c,-16'h007a,16'h0078,-16'h005d,-16'h0045,-16'h0014,16'h006d,-16'h0001,-16'h0009,16'h0000,16'h005c,-16'h001d,-16'h001a,-16'h002b,16'h0018,16'h0020,-16'h0025,16'h000e,16'h000f,-16'h0038,16'h0050,16'h001d,16'h005a,-16'h004a,-16'h000f,16'h0005,16'h0017,-16'h0083,16'h0007,16'h0037,16'h0002,-16'h000b,16'h0000,16'h0069,-16'h000a,-16'h0061,16'h0018,-16'h001f,16'h000e,16'h001c,-16'h0002,16'h0001,-16'h0021,-16'h0021,16'h0000,16'h0035,16'h0017,-16'h0004,-16'h0051,-16'h002f,16'h002d,16'h0024,-16'h0004,16'h0046,-16'h0022,-16'h0044,16'h005f,16'h0004,-16'h0021,-16'h0034,-16'h0033,16'h0035,16'h0039,-16'h003f,-16'h0046,-16'h007f,16'h0067,-16'h0030,-16'h0050,-16'h0001,16'h006e,-16'h000b,-16'h0018,-16'h0013,16'h0046,-16'h0030,-16'h0024,-16'h001b,16'h0015,16'h0038,-16'h0019,-16'h0005,16'h001e,-16'h0035,16'h004c,16'h0002,16'h006f,-16'h0052,-16'h002f,-16'h002f,-16'h0008,-16'h001d,16'h0024,16'h003a,16'h0012,-16'h0006,16'h0010,16'h005a,-16'h0007,-16'h0088,16'h0013,-16'h000c,-16'h0003,16'h0082,-16'h001d,-16'h0016,-16'h0036,-16'h0007,-16'h0012,16'h0036,-16'h0022,16'h001b,-16'h003a,-16'h0015,16'h0018,16'h0016,16'h0016,16'h0051,-16'h0018,-16'h002a,16'h0008,-16'h001d,-16'h002c,-16'h003a,-16'h0028,16'h002b,16'h0022,-16'h0024,-16'h004f,-16'h0090,16'h005a,-16'h003a,-16'h0043,16'h0003,16'h0043,-16'h003c,-16'h000a,-16'h0007,16'h004d,-16'h0019,-16'h0019,-16'h000e,-16'h000c,16'h0024,-16'h0012,-16'h002a,16'h001a,-16'h002e,16'h004f,16'h0003,16'h0063,-16'h0064,16'h0006,-16'h0035,-16'h0001,16'h0048,16'h0020,16'h003d,16'h0009,-16'h0011,16'h001d,16'h0040,-16'h0012,-16'h0055,-16'h002b,16'h0005,16'h0012,16'h00a2,16'h0003,-16'h0035,-16'h005e,16'h0042,-16'h0023,16'h003e,-16'h002c,16'h0007,16'h0008,-16'h0029,16'h0024,16'h001e,16'h0005,16'h0086,16'h0005,-16'h002d,16'h000a,-16'h0002,-16'h0028,-16'h0038,-16'h0044,16'h003b,16'h0025,-16'h0041,-16'h0044,-16'h0056,16'h0031,-16'h0011,-16'h0044,-16'h001d,16'h005c,-16'h0078,-16'h0011,16'h0007,16'h0048,-16'h0013,-16'h0015,-16'h0009,16'h0010,16'h0036,16'h000a,-16'h001f,16'h0016,-16'h0035,16'h000a,-16'h005c,16'h0040,-16'h0073,16'h0021,16'h0000,16'h0006,16'h005d,16'h0018,-16'h0002,-16'h0004,-16'h0009,16'h004c,16'h0023,-16'h000e,-16'h0007,-16'h005f,16'h0000,-16'h000e,16'h0082,16'h001e,-16'h004e,-16'h003e,16'h0027,-16'h0039,16'h0034,-16'h001b,16'h0007,16'h0019,-16'h003d,16'h0011,16'h0031,-16'h000e,16'h0088,-16'h0021,-16'h0016,16'h0005,-16'h0012,-16'h0019,-16'h006b,-16'h0037,16'h002c,16'h002b,-16'h0021,-16'h0030,-16'h0016,16'h0016,-16'h000a,-16'h0057,-16'h001f,16'h0070,-16'h0057,-16'h0027,-16'h0008,16'h003d,16'h000f,-16'h000e,16'h002d,-16'h000c,16'h002e,16'h0019,-16'h003d,16'h0013,-16'h0002,16'h0022,-16'h0057,16'h000e,-16'h007e,16'h0007,-16'h0012,16'h000b,16'h0071,-16'h0015,-16'h001e,-16'h0034,16'h0032,16'h0039,16'h0005,16'h0000,16'h003c,-16'h008d,16'h0019,-16'h0024,16'h0075,16'h001a,-16'h006e,-16'h0021,16'h006f,-16'h003e,16'h001f,-16'h0002,-16'h0014,16'h0021,-16'h0044,16'h0028,16'h000d,-16'h000d,16'h0093,-16'h0021,16'h0010,-16'h0056,-16'h0005,16'h0005,-16'h0045,-16'h007b,16'h0049,16'h0031,-16'h0012,-16'h002a,16'h000c,-16'h0027,16'h0008,-16'h0079,-16'h003e,16'h0048,-16'h0058,-16'h0037,16'h0000,16'h0054,16'h0000,-16'h0009,16'h0026,16'h000e,16'h0015,16'h002f,-16'h0022,-16'h001e,-16'h001e,16'h003d,-16'h003d,-16'h001f,-16'h009d,16'h003b,-16'h0013,-16'h0026,16'h003b,-16'h0018,-16'h0019,-16'h0037,16'h0024,16'h0038,-16'h003b,16'h001e,16'h007e,-16'h008e,16'h002b,-16'h0021,16'h007a,16'h002b,-16'h0042,16'h0000,16'h006a,-16'h005e,-16'h0007,16'h0027,16'h0000,16'h0057,-16'h0010,16'h0023,16'h001c,-16'h0010,16'h009a,-16'h001e,16'h0017,-16'h007a,16'h0007,16'h0001,-16'h003e,-16'h00a3,16'h0041,16'h0030,-16'h0005,-16'h004e,16'h001f,-16'h0008,16'h001b,-16'h00ac,-16'h002b,16'h0005,-16'h0065,-16'h004e,-16'h0009,16'h0032,16'h000f,16'h0001,16'h0023,16'h0004,16'h0003,16'h004a,-16'h0010,-16'h0017,16'h0006,16'h002a,-16'h0044,-16'h0016,-16'h0099,16'h0051,-16'h0013,-16'h0034,16'h003f,-16'h0048,-16'h0053,-16'h001c,16'h0013,16'h0037,-16'h0044,16'h002c,16'h0070,-16'h006d,16'h001b,-16'h0029,16'h0024,16'h002f,-16'h0031,16'h0056,16'h0058,-16'h002c,16'h0009,16'h0077,-16'h003c,16'h0057,-16'h0017,16'h001f,16'h0035,-16'h0005,16'h009d,-16'h0040,16'h0014,-16'h004b,16'h0000,-16'h000d,-16'h0044,-16'h00aa,16'h0054,16'h0039,-16'h002a,-16'h005c,16'h0038,16'h0021,-16'h0007,-16'h00af,-16'h001a,-16'h0021,-16'h0044,-16'h0043,16'h002e,16'h004a,16'h001a,16'h0036,16'h003e,16'h0017,16'h0016,16'h004e,16'h0001,16'h0005,16'h0021,16'h0025,-16'h0031,-16'h0027,-16'h0082,16'h005a,16'h001c,-16'h005a,16'h0037,-16'h0062,-16'h0036,-16'h0041,16'h000c,16'h000a,-16'h0020,16'h003c,16'h0033,-16'h0068,16'h000e,-16'h0008,-16'h001a,16'h002b,-16'h0017,16'h0050,16'h003d,-16'h0041,16'h0021,16'h007b,-16'h003d,16'h006e,-16'h001b,16'h0033,16'h001d,16'h0034,16'h008b,-16'h0006,16'h002d,-16'h0039,16'h0019,-16'h0021,-16'h002f,-16'h00b2,16'h0069,16'h0036,-16'h003f,-16'h0052,16'h0028,16'h0074,16'h000a,-16'h00ec,16'h0000,-16'h0023,-16'h000d,-16'h004c,-16'h000d,16'h0039,16'h0021,16'h004f,16'h0034,16'h000f,16'h0000,16'h005f,-16'h000b,-16'h000b,16'h000e,16'h001e,-16'h000d,-16'h0017,-16'h0088,16'h0046,-16'h0018,-16'h005b,16'h000e,-16'h0099,-16'h0043,-16'h002b,16'h000b,-16'h0003,-16'h004d,16'h0020,16'h0032,-16'h008c,16'h002f,-16'h002c,-16'h0054,16'h0021,16'h0003,16'h0042,16'h0064,-16'h0027,16'h0020,16'h0056,-16'h004b,-16'h000f,16'h001a,16'h002c,16'h0030,16'h0037,16'h006e,-16'h0009,16'h000c,-16'h0037,16'h0027,-16'h0013,16'h0005,-16'h0062,16'h006d,16'h0032,-16'h0044,-16'h006c,16'h002f,16'h005c,16'h002b,-16'h0105,-16'h0018,-16'h0036,16'h0016,-16'h001e,-16'h003f,16'h0017,-16'h0023,16'h0078,16'h0032,16'h003e,16'h0023,16'h0048,16'h0003,-16'h0029,-16'h001d,16'h001a,-16'h0021,16'h002b,-16'h0080,16'h005b,-16'h0030,-16'h0097,16'h0050,-16'h0090,-16'h0075,-16'h0031,16'h0001,-16'h003a,-16'h004d,16'h0034,16'h002d,-16'h003c,16'h0017,-16'h0017,-16'h0025,16'h001f,16'h000e,16'h0028,16'h0037,16'h0007,16'h0042,16'h000f,-16'h004b,-16'h0041,16'h003d,16'h004d,16'h0024,16'h0081,16'h0051,-16'h0004,-16'h0008,-16'h0058,16'h0011,-16'h0004,-16'h0007,-16'h0049,16'h0065,16'h0010,-16'h0058,-16'h005b,16'h001f,16'h0085,16'h0021,-16'h0112,-16'h002a,-16'h0059,-16'h000d,-16'h0019,-16'h003a,16'h002a,-16'h0049,16'h006b,16'h003a,16'h001f,16'h000c,16'h0028,16'h0000,-16'h0024,16'h0006,-16'h002f,-16'h0015,16'h003d,-16'h0093,16'h006c,-16'h001c,-16'h0099,16'h0053,-16'h00a4,-16'h0065,-16'h0042,16'h002d,-16'h0041,-16'h002d,16'h0019,16'h000c,-16'h0030,-16'h0020,-16'h0024,-16'h000d,16'h000c,16'h001b,16'h0005,16'h003f,16'h0028,16'h0065,16'h000a,16'h0016,-16'h0063,16'h0023,16'h007a,16'h0018,16'h007c,16'h003f,16'h0000,16'h000d,-16'h0039,16'h0018,-16'h0022,-16'h0020,-16'h002a,16'h0057,16'h0015,-16'h0047,-16'h0057,16'h000b,16'h00a1,16'h003c,-16'h0103,-16'h003f,-16'h006b,-16'h001d,16'h002e,-16'h0036,16'h0009,-16'h0091,16'h006a,16'h0050,16'h0014,16'h0006,16'h0003,-16'h000e,-16'h0023,-16'h0019,-16'h0037,16'h0003,16'h0047,-16'h0087,16'h006a,16'h0000,-16'h0084,16'h002a,-16'h00a7,-16'h004f,-16'h0041,16'h0060,-16'h0022,-16'h004e,16'h0027,-16'h000a,-16'h0030,-16'h00ba,16'h0010,16'h0005,16'h000a,-16'h001b,16'h0003,16'h0030,16'h0054,16'h0087,-16'h0009,16'h0012,-16'h004b,16'h0079,16'h0078,-16'h0006,16'h0081,16'h003a,-16'h0004,16'h0012,-16'h0041,16'h000b,-16'h0022,-16'h003e,-16'h0058,16'h0045,-16'h000f,-16'h0083,-16'h003d,16'h0017,16'h007b,16'h0014,-16'h0103,-16'h002a,-16'h00b8,-16'h001f,16'h0022,16'h0000,-16'h000a,-16'h0051,16'h005a,16'h0037,16'h0001,16'h0019,-16'h0017,-16'h000d,-16'h0030,-16'h0030,-16'h005e,16'h002d,16'h005a,-16'h0082,16'h0023,16'h0015,-16'h0080,16'h000e,-16'h009e,-16'h0036,-16'h004d,16'h0047,-16'h0029,-16'h0073,16'h0039,-16'h000c,-16'h0040,-16'h00fd,16'h0007,16'h001b,16'h001f,-16'h001b,-16'h000c,16'h003d,16'h0073,16'h0092,-16'h000d,16'h002a,-16'h0024,16'h007f,16'h007c,-16'h003a,16'h0078,16'h001a,-16'h0009,16'h0034,-16'h004c,16'h0023,16'h0003,-16'h0024,-16'h0044,16'h0051,-16'h0020,-16'h007e,-16'h001e,-16'h0001,16'h0024,16'h0011,-16'h00f1,-16'h0014,-16'h00cf,16'h0004,16'h0026,16'h0036,-16'h001e,-16'h0035,16'h0024,16'h0035,16'h000d,16'h0004,-16'h0036,16'h000d,-16'h0048,-16'h002a,-16'h0030,16'h0031,16'h003e,-16'h00a1,16'h001f,16'h0020,-16'h009d,-16'h0058,-16'h00a0,-16'h000c,-16'h005c,16'h0049,-16'h0003,-16'h0091,16'h004a,16'h0001,-16'h0052,-16'h00ce,16'h0015,16'h0037,16'h0010,-16'h0029,16'h000f,16'h004b,16'h0082,16'h009c,-16'h0010,16'h0042,16'h0030,16'h007c,16'h00bb,-16'h0035,16'h0062,-16'h0006,-16'h000b,16'h001e,-16'h0039,16'h0021,16'h000f,-16'h001c,-16'h002d,16'h0049,16'h0000,-16'h008f,-16'h0017,-16'h0003,-16'h0004,-16'h0025,-16'h00da,16'h0005,-16'h00b8,16'h001f,16'h0058,16'h0019,-16'h0042,-16'h0005,16'h0015,16'h0021,16'h0005,16'h0026,-16'h0030,16'h001e,-16'h003c,-16'h0008,-16'h0014,16'h004b,16'h0035,-16'h0094,16'h003f,16'h000d,-16'h0064,-16'h0033,-16'h0084,16'h0020,-16'h0041,16'h0052,16'h0008,-16'h007d,16'h0062,-16'h0024,-16'h005e,-16'h005b,-16'h000f,16'h0037,-16'h0040,-16'h000e,-16'h001c,16'h0047,16'h0068,16'h00ac,16'h0009,16'h005b,16'h0054,16'h004c,16'h00c2,-16'h005e,16'h0058,16'h0008,-16'h0008,16'h0015,-16'h0027,16'h0007,16'h0024,-16'h0024,16'h003f,16'h0059,-16'h0029,-16'h0064,-16'h0014,16'h000f,-16'h0027,-16'h0045,-16'h009f,16'h0017,-16'h0078,16'h002d,16'h0035,16'h0034,-16'h0062,-16'h0015,16'h0019,16'h001e,16'h0025,16'h0034,-16'h0025,16'h0051,-16'h003b,-16'h0017,-16'h0015,16'h0075,16'h002a,-16'h0079,16'h0021,16'h000e,-16'h0030,-16'h0027,-16'h0074,16'h0017,-16'h0020,16'h003c,16'h0014,-16'h0064,16'h0060,-16'h0043,-16'h0044,-16'h0041,16'h0001,-16'h0001,-16'h007a,-16'h0010,-16'h002e,16'h0043,16'h006b,16'h005a,16'h0007,16'h002e,16'h0020,16'h004e,16'h00ba,-16'h008c,16'h004a,16'h000d,-16'h001c,16'h000d,-16'h0032,16'h0010,16'h003a,-16'h001b,16'h0068,16'h0033,-16'h0029,-16'h0056,-16'h0017,16'h0023,-16'h003e,-16'h005e,-16'h00aa,16'h0005,-16'h0035,16'h0025,16'h0024,16'h002a,-16'h0069,-16'h0011,-16'h0004,16'h0007,16'h002c,16'h002b,-16'h0027,16'h0033,-16'h0016,-16'h0006,-16'h0016,16'h00a1,16'h0033,-16'h0089,16'h001f,16'h0017,-16'h0022,16'h0010,-16'h004f,16'h0023,-16'h0018,16'h003d,16'h0038,-16'h004c,16'h003c,-16'h004c,-16'h0021,-16'h0009,16'h0004,16'h0019,-16'h005e,-16'h000c,-16'h0048,16'h001f,16'h001e,16'h0054,16'h0025,16'h0017,16'h0038,16'h000e,16'h008b,-16'h0066,16'h0043,-16'h0003,-16'h0011,-16'h0012,-16'h000f,16'h000a,16'h002f,-16'h0032,16'h0075,16'h0018,-16'h002d,-16'h0048,-16'h0002,16'h005e,-16'h0010,-16'h004d,-16'h007b,-16'h000f,-16'h0018,16'h002d,16'h0039,16'h0021,-16'h0034,16'h000a,16'h0000,16'h000f,16'h001b,16'h0021,-16'h0009,16'h005a,-16'h000f,-16'h000c,-16'h002f,16'h0093,16'h0000,-16'h0082,16'h001e,16'h0000,-16'h000b,16'h0017,-16'h0039,16'h0023,16'h000b,16'h0029,16'h002d,-16'h0022,16'h0036,-16'h0031,-16'h0008,-16'h0005,16'h0013,-16'h0002,-16'h0055,-16'h000c,-16'h0030,-16'h0002,16'h0013,16'h000c,16'h001a,-16'h0001,16'h0027,-16'h0021,16'h007c,-16'h0059,16'h005b,16'h0001,16'h0002,-16'h0006,-16'h0002,16'h0020,-16'h0019,-16'h0010,16'h0073,16'h000f,-16'h0005,-16'h001d,16'h0005,16'h007c,-16'h001b,-16'h0044,-16'h0059,-16'h0006,-16'h0016,-16'h0001,16'h0018,16'h000e,-16'h001e,16'h001a,16'h0010,16'h0023,16'h000d,16'h0004,16'h000f,16'h005a,16'h0007,16'h0011,-16'h0007,16'h006e,16'h0023,-16'h0061,-16'h000d,-16'h0007,-16'h0006,16'h0012,-16'h0004,16'h0027,16'h0004,16'h000b,16'h0018,16'h0003,16'h0000,-16'h002f,-16'h0016,16'h0003,16'h001f,-16'h0017,-16'h002f,16'h0010,-16'h0017,-16'h0010,-16'h000e,16'h0015,16'h001d,16'h0000,-16'h0009,-16'h0024,16'h0061,-16'h002b,16'h005a,-16'h0006,-16'h0003,-16'h001d,-16'h0002,16'h0013,16'h0009,-16'h0027,16'h003f,16'h0017,-16'h0007,-16'h0019,16'h0002,16'h0053,-16'h0017,-16'h002c,-16'h0047,16'h0019,16'h000d,-16'h000a,16'h000b};
    localparam [1023:0] bias_0 = {16'h0077,-16'h00d9,-16'h001a,-16'h003b,-16'h003f,16'h0098,16'h0006,-16'h00a6,-16'h01d4,-16'h0145,16'h0051,16'h00ce,-16'h00df,16'h000a,-16'h001a,16'h007e,16'h00d5,-16'h014e,16'h011a,-16'h0018,16'h0150,-16'h01f4,-16'h0064,-16'h0013,16'h002b,-16'h00b5,16'h001d,16'h0000,16'h002f,-16'h002f,16'h0115,16'h000d,-16'h00c3,16'h00bf,-16'h0030,16'h00e9,16'h0078,16'h00c5,-16'h0194,16'h006f,16'h005f,-16'h00ef,-16'h007d,-16'h0106,16'h001c,-16'h0029,-16'h008e,16'h0062,-16'h0119,16'h009c,-16'h0039,-16'h0102,-16'h01cb,16'h0074,16'h0072,-16'h00f5,-16'h00f0,-16'h0071,-16'h016d,-16'h00a6,-16'h0180,-16'h010c,16'h0040,-16'h004b};

    localparam SWAIT = 3'd0;
    localparam SDOT = 3'd1;
    localparam SBIAS = 3'd2;
    localparam SRELU = 3'd3;
    localparam SFIN = 3'd4;
    reg [2:0] state, next_state;

    reg  [16 - 1:0]     row, next_row;
    reg  [16*64 - 1:0]  next_layer_0;
    reg                 next_finish;
    wire [16 - 1:0]     curr_input_digit;

    assign curr_input_digit = {15'b0,layer_input[row]};
    /* ------------------------------------Sequential------------------------------------- */
    always @(posedge clk ) begin
        if(rst) begin
            state <= SWAIT;
            row <= 0;
            layer_0 <= 0;
            finish <= 0;
        end else begin
            state <= next_state;
            row <= next_row;
            layer_0 <= next_layer_0;
            finish <= next_finish;
        end
    end
    /* ------------------------------------State Combinational------------------------------------- */
    always @(*) begin
        case (state)
            SWAIT: begin
                if(start) next_state = SDOT;
                else next_state = state;
            end
            SDOT: begin
                if(row == HEIGHT - 1) next_state = SBIAS;
                else next_state = state;
            end
            SBIAS: next_state = SRELU;
            SRELU: next_state = SFIN;
            default: next_state = SWAIT;
        endcase
    end
    /* ------------------------------------Other Combinationals------------------------------------- */
    always @(*) begin
        case (state)
            SDOT: next_row = row + 16'b1;
            default: next_row = 16'b0;
        endcase
    end
    // finish
    always @(*) begin
        case (state)
            SRELU: next_finish = 1'b1;
            default: next_finish = 1'b0;
        endcase
    end
    /* ------------------------------------Layer Calculation------------------------------------- */
    always @(*) begin
        case (state)
            SWAIT: begin
                if(start) next_layer_0 = 0;
                else next_layer_0 = layer_0;
            end
            SDOT: begin
                next_layer_0[15-:16] = layer_0[15-:16] + (curr_input_digit * kernel_0[(row*64+0+1)*16-1-:16]);
                next_layer_0[31-:16] = layer_0[31-:16] + (curr_input_digit * kernel_0[(row*64+1+1)*16-1-:16]);
                next_layer_0[47-:16] = layer_0[47-:16] + (curr_input_digit * kernel_0[(row*64+2+1)*16-1-:16]);
                next_layer_0[63-:16] = layer_0[63-:16] + (curr_input_digit * kernel_0[(row*64+3+1)*16-1-:16]);
                next_layer_0[79-:16] = layer_0[79-:16] + (curr_input_digit * kernel_0[(row*64+4+1)*16-1-:16]);
                next_layer_0[95-:16] = layer_0[95-:16] + (curr_input_digit * kernel_0[(row*64+5+1)*16-1-:16]);
                next_layer_0[111-:16] = layer_0[111-:16] + (curr_input_digit * kernel_0[(row*64+6+1)*16-1-:16]);
                next_layer_0[127-:16] = layer_0[127-:16] + (curr_input_digit * kernel_0[(row*64+7+1)*16-1-:16]);
                next_layer_0[143-:16] = layer_0[143-:16] + (curr_input_digit * kernel_0[(row*64+8+1)*16-1-:16]);
                next_layer_0[159-:16] = layer_0[159-:16] + (curr_input_digit * kernel_0[(row*64+9+1)*16-1-:16]);
                next_layer_0[175-:16] = layer_0[175-:16] + (curr_input_digit * kernel_0[(row*64+10+1)*16-1-:16]);
                next_layer_0[191-:16] = layer_0[191-:16] + (curr_input_digit * kernel_0[(row*64+11+1)*16-1-:16]);
                next_layer_0[207-:16] = layer_0[207-:16] + (curr_input_digit * kernel_0[(row*64+12+1)*16-1-:16]);
                next_layer_0[223-:16] = layer_0[223-:16] + (curr_input_digit * kernel_0[(row*64+13+1)*16-1-:16]);
                next_layer_0[239-:16] = layer_0[239-:16] + (curr_input_digit * kernel_0[(row*64+14+1)*16-1-:16]);
                next_layer_0[255-:16] = layer_0[255-:16] + (curr_input_digit * kernel_0[(row*64+15+1)*16-1-:16]);
                next_layer_0[271-:16] = layer_0[271-:16] + (curr_input_digit * kernel_0[(row*64+16+1)*16-1-:16]);
                next_layer_0[287-:16] = layer_0[287-:16] + (curr_input_digit * kernel_0[(row*64+17+1)*16-1-:16]);
                next_layer_0[303-:16] = layer_0[303-:16] + (curr_input_digit * kernel_0[(row*64+18+1)*16-1-:16]);
                next_layer_0[319-:16] = layer_0[319-:16] + (curr_input_digit * kernel_0[(row*64+19+1)*16-1-:16]);
                next_layer_0[335-:16] = layer_0[335-:16] + (curr_input_digit * kernel_0[(row*64+20+1)*16-1-:16]);
                next_layer_0[351-:16] = layer_0[351-:16] + (curr_input_digit * kernel_0[(row*64+21+1)*16-1-:16]);
                next_layer_0[367-:16] = layer_0[367-:16] + (curr_input_digit * kernel_0[(row*64+22+1)*16-1-:16]);
                next_layer_0[383-:16] = layer_0[383-:16] + (curr_input_digit * kernel_0[(row*64+23+1)*16-1-:16]);
                next_layer_0[399-:16] = layer_0[399-:16] + (curr_input_digit * kernel_0[(row*64+24+1)*16-1-:16]);
                next_layer_0[415-:16] = layer_0[415-:16] + (curr_input_digit * kernel_0[(row*64+25+1)*16-1-:16]);
                next_layer_0[431-:16] = layer_0[431-:16] + (curr_input_digit * kernel_0[(row*64+26+1)*16-1-:16]);
                next_layer_0[447-:16] = layer_0[447-:16] + (curr_input_digit * kernel_0[(row*64+27+1)*16-1-:16]);
                next_layer_0[463-:16] = layer_0[463-:16] + (curr_input_digit * kernel_0[(row*64+28+1)*16-1-:16]);
                next_layer_0[479-:16] = layer_0[479-:16] + (curr_input_digit * kernel_0[(row*64+29+1)*16-1-:16]);
                next_layer_0[495-:16] = layer_0[495-:16] + (curr_input_digit * kernel_0[(row*64+30+1)*16-1-:16]);
                next_layer_0[511-:16] = layer_0[511-:16] + (curr_input_digit * kernel_0[(row*64+31+1)*16-1-:16]);
                next_layer_0[527-:16] = layer_0[527-:16] + (curr_input_digit * kernel_0[(row*64+32+1)*16-1-:16]);
                next_layer_0[543-:16] = layer_0[543-:16] + (curr_input_digit * kernel_0[(row*64+33+1)*16-1-:16]);
                next_layer_0[559-:16] = layer_0[559-:16] + (curr_input_digit * kernel_0[(row*64+34+1)*16-1-:16]);
                next_layer_0[575-:16] = layer_0[575-:16] + (curr_input_digit * kernel_0[(row*64+35+1)*16-1-:16]);
                next_layer_0[591-:16] = layer_0[591-:16] + (curr_input_digit * kernel_0[(row*64+36+1)*16-1-:16]);
                next_layer_0[607-:16] = layer_0[607-:16] + (curr_input_digit * kernel_0[(row*64+37+1)*16-1-:16]);
                next_layer_0[623-:16] = layer_0[623-:16] + (curr_input_digit * kernel_0[(row*64+38+1)*16-1-:16]);
                next_layer_0[639-:16] = layer_0[639-:16] + (curr_input_digit * kernel_0[(row*64+39+1)*16-1-:16]);
                next_layer_0[655-:16] = layer_0[655-:16] + (curr_input_digit * kernel_0[(row*64+40+1)*16-1-:16]);
                next_layer_0[671-:16] = layer_0[671-:16] + (curr_input_digit * kernel_0[(row*64+41+1)*16-1-:16]);
                next_layer_0[687-:16] = layer_0[687-:16] + (curr_input_digit * kernel_0[(row*64+42+1)*16-1-:16]);
                next_layer_0[703-:16] = layer_0[703-:16] + (curr_input_digit * kernel_0[(row*64+43+1)*16-1-:16]);
                next_layer_0[719-:16] = layer_0[719-:16] + (curr_input_digit * kernel_0[(row*64+44+1)*16-1-:16]);
                next_layer_0[735-:16] = layer_0[735-:16] + (curr_input_digit * kernel_0[(row*64+45+1)*16-1-:16]);
                next_layer_0[751-:16] = layer_0[751-:16] + (curr_input_digit * kernel_0[(row*64+46+1)*16-1-:16]);
                next_layer_0[767-:16] = layer_0[767-:16] + (curr_input_digit * kernel_0[(row*64+47+1)*16-1-:16]);
                next_layer_0[783-:16] = layer_0[783-:16] + (curr_input_digit * kernel_0[(row*64+48+1)*16-1-:16]);
                next_layer_0[799-:16] = layer_0[799-:16] + (curr_input_digit * kernel_0[(row*64+49+1)*16-1-:16]);
                next_layer_0[815-:16] = layer_0[815-:16] + (curr_input_digit * kernel_0[(row*64+50+1)*16-1-:16]);
                next_layer_0[831-:16] = layer_0[831-:16] + (curr_input_digit * kernel_0[(row*64+51+1)*16-1-:16]);
                next_layer_0[847-:16] = layer_0[847-:16] + (curr_input_digit * kernel_0[(row*64+52+1)*16-1-:16]);
                next_layer_0[863-:16] = layer_0[863-:16] + (curr_input_digit * kernel_0[(row*64+53+1)*16-1-:16]);
                next_layer_0[879-:16] = layer_0[879-:16] + (curr_input_digit * kernel_0[(row*64+54+1)*16-1-:16]);
                next_layer_0[895-:16] = layer_0[895-:16] + (curr_input_digit * kernel_0[(row*64+55+1)*16-1-:16]);
                next_layer_0[911-:16] = layer_0[911-:16] + (curr_input_digit * kernel_0[(row*64+56+1)*16-1-:16]);
                next_layer_0[927-:16] = layer_0[927-:16] + (curr_input_digit * kernel_0[(row*64+57+1)*16-1-:16]);
                next_layer_0[943-:16] = layer_0[943-:16] + (curr_input_digit * kernel_0[(row*64+58+1)*16-1-:16]);
                next_layer_0[959-:16] = layer_0[959-:16] + (curr_input_digit * kernel_0[(row*64+59+1)*16-1-:16]);
                next_layer_0[975-:16] = layer_0[975-:16] + (curr_input_digit * kernel_0[(row*64+60+1)*16-1-:16]);
                next_layer_0[991-:16] = layer_0[991-:16] + (curr_input_digit * kernel_0[(row*64+61+1)*16-1-:16]);
                next_layer_0[1007-:16] = layer_0[1007-:16] + (curr_input_digit * kernel_0[(row*64+62+1)*16-1-:16]);
                next_layer_0[1023-:16] = layer_0[1023-:16] + (curr_input_digit * kernel_0[(row*64+63+1)*16-1-:16]);
            end
            SBIAS: begin
                next_layer_0[15-:16] = layer_0[15-:16] + bias_0[15-:16];
                next_layer_0[31-:16] = layer_0[31-:16] + bias_0[31-:16];
                next_layer_0[47-:16] = layer_0[47-:16] + bias_0[47-:16];
                next_layer_0[63-:16] = layer_0[63-:16] + bias_0[63-:16];
                next_layer_0[79-:16] = layer_0[79-:16] + bias_0[79-:16];
                next_layer_0[95-:16] = layer_0[95-:16] + bias_0[95-:16];
                next_layer_0[111-:16] = layer_0[111-:16] + bias_0[111-:16];
                next_layer_0[127-:16] = layer_0[127-:16] + bias_0[127-:16];
                next_layer_0[143-:16] = layer_0[143-:16] + bias_0[143-:16];
                next_layer_0[159-:16] = layer_0[159-:16] + bias_0[159-:16];
                next_layer_0[175-:16] = layer_0[175-:16] + bias_0[175-:16];
                next_layer_0[191-:16] = layer_0[191-:16] + bias_0[191-:16];
                next_layer_0[207-:16] = layer_0[207-:16] + bias_0[207-:16];
                next_layer_0[223-:16] = layer_0[223-:16] + bias_0[223-:16];
                next_layer_0[239-:16] = layer_0[239-:16] + bias_0[239-:16];
                next_layer_0[255-:16] = layer_0[255-:16] + bias_0[255-:16];
                next_layer_0[271-:16] = layer_0[271-:16] + bias_0[271-:16];
                next_layer_0[287-:16] = layer_0[287-:16] + bias_0[287-:16];
                next_layer_0[303-:16] = layer_0[303-:16] + bias_0[303-:16];
                next_layer_0[319-:16] = layer_0[319-:16] + bias_0[319-:16];
                next_layer_0[335-:16] = layer_0[335-:16] + bias_0[335-:16];
                next_layer_0[351-:16] = layer_0[351-:16] + bias_0[351-:16];
                next_layer_0[367-:16] = layer_0[367-:16] + bias_0[367-:16];
                next_layer_0[383-:16] = layer_0[383-:16] + bias_0[383-:16];
                next_layer_0[399-:16] = layer_0[399-:16] + bias_0[399-:16];
                next_layer_0[415-:16] = layer_0[415-:16] + bias_0[415-:16];
                next_layer_0[431-:16] = layer_0[431-:16] + bias_0[431-:16];
                next_layer_0[447-:16] = layer_0[447-:16] + bias_0[447-:16];
                next_layer_0[463-:16] = layer_0[463-:16] + bias_0[463-:16];
                next_layer_0[479-:16] = layer_0[479-:16] + bias_0[479-:16];
                next_layer_0[495-:16] = layer_0[495-:16] + bias_0[495-:16];
                next_layer_0[511-:16] = layer_0[511-:16] + bias_0[511-:16];
                next_layer_0[527-:16] = layer_0[527-:16] + bias_0[527-:16];
                next_layer_0[543-:16] = layer_0[543-:16] + bias_0[543-:16];
                next_layer_0[559-:16] = layer_0[559-:16] + bias_0[559-:16];
                next_layer_0[575-:16] = layer_0[575-:16] + bias_0[575-:16];
                next_layer_0[591-:16] = layer_0[591-:16] + bias_0[591-:16];
                next_layer_0[607-:16] = layer_0[607-:16] + bias_0[607-:16];
                next_layer_0[623-:16] = layer_0[623-:16] + bias_0[623-:16];
                next_layer_0[639-:16] = layer_0[639-:16] + bias_0[639-:16];
                next_layer_0[655-:16] = layer_0[655-:16] + bias_0[655-:16];
                next_layer_0[671-:16] = layer_0[671-:16] + bias_0[671-:16];
                next_layer_0[687-:16] = layer_0[687-:16] + bias_0[687-:16];
                next_layer_0[703-:16] = layer_0[703-:16] + bias_0[703-:16];
                next_layer_0[719-:16] = layer_0[719-:16] + bias_0[719-:16];
                next_layer_0[735-:16] = layer_0[735-:16] + bias_0[735-:16];
                next_layer_0[751-:16] = layer_0[751-:16] + bias_0[751-:16];
                next_layer_0[767-:16] = layer_0[767-:16] + bias_0[767-:16];
                next_layer_0[783-:16] = layer_0[783-:16] + bias_0[783-:16];
                next_layer_0[799-:16] = layer_0[799-:16] + bias_0[799-:16];
                next_layer_0[815-:16] = layer_0[815-:16] + bias_0[815-:16];
                next_layer_0[831-:16] = layer_0[831-:16] + bias_0[831-:16];
                next_layer_0[847-:16] = layer_0[847-:16] + bias_0[847-:16];
                next_layer_0[863-:16] = layer_0[863-:16] + bias_0[863-:16];
                next_layer_0[879-:16] = layer_0[879-:16] + bias_0[879-:16];
                next_layer_0[895-:16] = layer_0[895-:16] + bias_0[895-:16];
                next_layer_0[911-:16] = layer_0[911-:16] + bias_0[911-:16];
                next_layer_0[927-:16] = layer_0[927-:16] + bias_0[927-:16];
                next_layer_0[943-:16] = layer_0[943-:16] + bias_0[943-:16];
                next_layer_0[959-:16] = layer_0[959-:16] + bias_0[959-:16];
                next_layer_0[975-:16] = layer_0[975-:16] + bias_0[975-:16];
                next_layer_0[991-:16] = layer_0[991-:16] + bias_0[991-:16];
                next_layer_0[1007-:16] = layer_0[1007-:16] + bias_0[1007-:16];
                next_layer_0[1023-:16] = layer_0[1023-:16] + bias_0[1023-:16];
            end
            SRELU: begin
                next_layer_0[15-:16] = (layer_0[15] ? 16'b0 : layer_0[15-:16]);
                next_layer_0[31-:16] = (layer_0[31] ? 16'b0 : layer_0[31-:16]);
                next_layer_0[47-:16] = (layer_0[47] ? 16'b0 : layer_0[47-:16]);
                next_layer_0[63-:16] = (layer_0[63] ? 16'b0 : layer_0[63-:16]);
                next_layer_0[79-:16] = (layer_0[79] ? 16'b0 : layer_0[79-:16]);
                next_layer_0[95-:16] = (layer_0[95] ? 16'b0 : layer_0[95-:16]);
                next_layer_0[111-:16] = (layer_0[111] ? 16'b0 : layer_0[111-:16]);
                next_layer_0[127-:16] = (layer_0[127] ? 16'b0 : layer_0[127-:16]);
                next_layer_0[143-:16] = (layer_0[143] ? 16'b0 : layer_0[143-:16]);
                next_layer_0[159-:16] = (layer_0[159] ? 16'b0 : layer_0[159-:16]);
                next_layer_0[175-:16] = (layer_0[175] ? 16'b0 : layer_0[175-:16]);
                next_layer_0[191-:16] = (layer_0[191] ? 16'b0 : layer_0[191-:16]);
                next_layer_0[207-:16] = (layer_0[207] ? 16'b0 : layer_0[207-:16]);
                next_layer_0[223-:16] = (layer_0[223] ? 16'b0 : layer_0[223-:16]);
                next_layer_0[239-:16] = (layer_0[239] ? 16'b0 : layer_0[239-:16]);
                next_layer_0[255-:16] = (layer_0[255] ? 16'b0 : layer_0[255-:16]);
                next_layer_0[271-:16] = (layer_0[271] ? 16'b0 : layer_0[271-:16]);
                next_layer_0[287-:16] = (layer_0[287] ? 16'b0 : layer_0[287-:16]);
                next_layer_0[303-:16] = (layer_0[303] ? 16'b0 : layer_0[303-:16]);
                next_layer_0[319-:16] = (layer_0[319] ? 16'b0 : layer_0[319-:16]);
                next_layer_0[335-:16] = (layer_0[335] ? 16'b0 : layer_0[335-:16]);
                next_layer_0[351-:16] = (layer_0[351] ? 16'b0 : layer_0[351-:16]);
                next_layer_0[367-:16] = (layer_0[367] ? 16'b0 : layer_0[367-:16]);
                next_layer_0[383-:16] = (layer_0[383] ? 16'b0 : layer_0[383-:16]);
                next_layer_0[399-:16] = (layer_0[399] ? 16'b0 : layer_0[399-:16]);
                next_layer_0[415-:16] = (layer_0[415] ? 16'b0 : layer_0[415-:16]);
                next_layer_0[431-:16] = (layer_0[431] ? 16'b0 : layer_0[431-:16]);
                next_layer_0[447-:16] = (layer_0[447] ? 16'b0 : layer_0[447-:16]);
                next_layer_0[463-:16] = (layer_0[463] ? 16'b0 : layer_0[463-:16]);
                next_layer_0[479-:16] = (layer_0[479] ? 16'b0 : layer_0[479-:16]);
                next_layer_0[495-:16] = (layer_0[495] ? 16'b0 : layer_0[495-:16]);
                next_layer_0[511-:16] = (layer_0[511] ? 16'b0 : layer_0[511-:16]);
                next_layer_0[527-:16] = (layer_0[527] ? 16'b0 : layer_0[527-:16]);
                next_layer_0[543-:16] = (layer_0[543] ? 16'b0 : layer_0[543-:16]);
                next_layer_0[559-:16] = (layer_0[559] ? 16'b0 : layer_0[559-:16]);
                next_layer_0[575-:16] = (layer_0[575] ? 16'b0 : layer_0[575-:16]);
                next_layer_0[591-:16] = (layer_0[591] ? 16'b0 : layer_0[591-:16]);
                next_layer_0[607-:16] = (layer_0[607] ? 16'b0 : layer_0[607-:16]);
                next_layer_0[623-:16] = (layer_0[623] ? 16'b0 : layer_0[623-:16]);
                next_layer_0[639-:16] = (layer_0[639] ? 16'b0 : layer_0[639-:16]);
                next_layer_0[655-:16] = (layer_0[655] ? 16'b0 : layer_0[655-:16]);
                next_layer_0[671-:16] = (layer_0[671] ? 16'b0 : layer_0[671-:16]);
                next_layer_0[687-:16] = (layer_0[687] ? 16'b0 : layer_0[687-:16]);
                next_layer_0[703-:16] = (layer_0[703] ? 16'b0 : layer_0[703-:16]);
                next_layer_0[719-:16] = (layer_0[719] ? 16'b0 : layer_0[719-:16]);
                next_layer_0[735-:16] = (layer_0[735] ? 16'b0 : layer_0[735-:16]);
                next_layer_0[751-:16] = (layer_0[751] ? 16'b0 : layer_0[751-:16]);
                next_layer_0[767-:16] = (layer_0[767] ? 16'b0 : layer_0[767-:16]);
                next_layer_0[783-:16] = (layer_0[783] ? 16'b0 : layer_0[783-:16]);
                next_layer_0[799-:16] = (layer_0[799] ? 16'b0 : layer_0[799-:16]);
                next_layer_0[815-:16] = (layer_0[815] ? 16'b0 : layer_0[815-:16]);
                next_layer_0[831-:16] = (layer_0[831] ? 16'b0 : layer_0[831-:16]);
                next_layer_0[847-:16] = (layer_0[847] ? 16'b0 : layer_0[847-:16]);
                next_layer_0[863-:16] = (layer_0[863] ? 16'b0 : layer_0[863-:16]);
                next_layer_0[879-:16] = (layer_0[879] ? 16'b0 : layer_0[879-:16]);
                next_layer_0[895-:16] = (layer_0[895] ? 16'b0 : layer_0[895-:16]);
                next_layer_0[911-:16] = (layer_0[911] ? 16'b0 : layer_0[911-:16]);
                next_layer_0[927-:16] = (layer_0[927] ? 16'b0 : layer_0[927-:16]);
                next_layer_0[943-:16] = (layer_0[943] ? 16'b0 : layer_0[943-:16]);
                next_layer_0[959-:16] = (layer_0[959] ? 16'b0 : layer_0[959-:16]);
                next_layer_0[975-:16] = (layer_0[975] ? 16'b0 : layer_0[975-:16]);
                next_layer_0[991-:16] = (layer_0[991] ? 16'b0 : layer_0[991-:16]);
                next_layer_0[1007-:16] = (layer_0[1007] ? 16'b0 : layer_0[1007-:16]);
                next_layer_0[1023-:16] = (layer_0[1023] ? 16'b0 : layer_0[1023-:16]);
            end
            SFIN: next_layer_0 = layer_0;
            default: next_layer_0 = layer_0;
        endcase
    end
endmodule