`timescale 1ps/1ps
module SudokuGenerator #(
    parameter size = 9,
    parameter bit = 4
    ) (
    input [15:0] random,
    output reg [81*4-1:0] board,
    output wire [81-1:0]  board_blank
    );
    
    genvar i;
    generate
        for(i = 0; i < 81; i = i + 1) begin
            assign board_blank[i] = board[(i+1)*bit-1-:bit] == 4'd0;
        end
    endgenerate

    always @(*) begin
        case (random[5:0])
            8'h00:board={4'd8,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd7,4'd7,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0};
            8'h01:board={4'd3,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd4,4'd9,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2};
            8'h02:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd2,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd9,4'd2,4'd3,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd4,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0};
            8'h03:board={4'd2,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd4,4'd0,4'd9,4'd0,4'd5,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd3,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0};
            8'h04:board={4'd0,4'd9,4'd0,4'd2,4'd0,4'd4,4'd5,4'd0,4'd0,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd9,4'd5,4'd0,4'd0,4'd8,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd9};
            8'h05:board={4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd6,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h06:board={4'd6,4'd1,4'd0,4'd8,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd6,4'd4,4'd0};
            8'h07:board={4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd2,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h08:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd2,4'd1,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0};
            8'h09:board={4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0};
            8'h0a:board={4'd1,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd0,4'd5,4'd3,4'd0,4'd0,4'd4,4'd3,4'd0,4'd5,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd5,4'd8,4'd0,4'd7,4'd0,4'd0};
            8'h0b:board={4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd8,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd6,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h0c:board={4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd8,4'd5,4'd0,4'd1,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3};
            8'h0d:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd5,4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0};
            8'h0e:board={4'd0,4'd0,4'd2,4'd0,4'd4,4'd5,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd6,4'd1,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0};
            8'h0f:board={4'd0,4'd0,4'd7,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd2,4'd4,4'd0,4'd6,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0};
            8'h10:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd3,4'd6,4'd1,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0};
            8'h11:board={4'd0,4'd6,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd2,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd7,4'd8};
            8'h12:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd1,4'd0,4'd9,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd5,4'd8,4'd0,4'd0,4'd0};
            8'h13:board={4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd9,4'd7,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0};
            8'h14:board={4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd1};
            8'h15:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0};
            8'h16:board={4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd4,4'd9,4'd0,4'd7,4'd5,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0};
            8'h17:board={4'd0,4'd3,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd1,4'd0,4'd2,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd7,4'd8,4'd0,4'd8,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd4,4'd1,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h18:board={4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd4,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd6,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd4,4'd0,4'd0};
            8'h19:board={4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd9,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3};
            8'h1a:board={4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd2,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd6,4'd2,4'd0,4'd0};
            8'h1b:board={4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd1,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd2,4'd5,4'd0,4'd7,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h1c:board={4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h1d:board={4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd9,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4};
            8'h1e:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd4,4'd3,4'd6,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd4,4'd0};
            8'h1f:board={4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd1,4'd0,4'd7,4'd8,4'd0,4'd2,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd6,4'd8,4'd5,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h20:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd2,4'd5,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd7,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0};
            8'h21:board={4'd8,4'd7,4'd0,4'd0,4'd0,4'd1,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd5,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9};
            8'h22:board={4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd3,4'd5,4'd0,4'd4,4'd6,4'd0,4'd9,4'd4,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3};
            8'h23:board={4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd5,4'd0,4'd6,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd1,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd7,4'd6};
            8'h24:board={4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd8,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h25:board={4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd7,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h26:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0};
            8'h27:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd8,4'd4,4'd3,4'd1,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0};
            8'h28:board={4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd5,4'd0,4'd0,4'd8,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd2,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0};
            8'h29:board={4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9};
            8'h2a:board={4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd1,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7,4'd3,4'd0,4'd0};
            8'h2b:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd9,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd8,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0};
            8'h2c:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd6,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3,4'd8,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd4,4'd9,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0};
            8'h2d:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd8,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5};
            8'h2e:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd8,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd8,4'd4,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd3};
            8'h2f:board={4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd7,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd6,4'd0,4'd1,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0};
            8'h30:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd4,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd9,4'd1,4'd8,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0};
            8'h31:board={4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd4,4'd2,4'd0,4'd9,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd4};
            8'h32:board={4'd4,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd2,4'd9,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4};
            8'h33:board={4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd5,4'd7,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd4,4'd8,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd3,4'd0};
            8'h34:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd5,4'd6,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd6,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0};
            8'h35:board={4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h36:board={4'd0,4'd1,4'd3,4'd4,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3};
            8'h37:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd3,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd7,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd9,4'd4,4'd0};
            8'h38:board={4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd3,4'd0,4'd8,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0};
            8'h39:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd6,4'd3,4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0};
            8'h3a:board={4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd8,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'h3b:board={4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd3,4'd1,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'h3c:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd3,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd1,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd2,4'd0,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h3d:board={4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd7,4'd0,4'd0,4'd4,4'd2,4'd6,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd5,4'd0,4'd4,4'd7,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h3e:board={4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd4,4'd0,4'd2,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd2,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd8,4'd0};
            8'h3f:board={4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0};
        endcase
    end
endmodule