`timescale 1ps/1ps
module Dense_1 (
    input a
    );
    
endmodule