`timescale 1ps/1ps
module SudokuGenerator #(
    parameter size = 9,
    parameter bit = 4
    ) (
    input [15:0] random,
    output reg [81*4-1:0] board
    );
    
    // localparam EASY = 2'd0;
    // localparam NORM = 2'd1;
    // localparam HARD = 2'd2;

    always @(*) begin
        case (random[7:0])
            8'h00:board={4'd8,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd7,4'd7,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0};
            8'h01:board={4'd3,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd4,4'd9,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2};
            8'h02:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd2,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd9,4'd2,4'd3,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd4,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0};
            8'h03:board={4'd2,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd4,4'd0,4'd9,4'd0,4'd5,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd3,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0};
            8'h04:board={4'd0,4'd9,4'd0,4'd2,4'd0,4'd4,4'd5,4'd0,4'd0,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd9,4'd5,4'd0,4'd0,4'd8,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd9};
            8'h05:board={4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd6,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h06:board={4'd6,4'd1,4'd0,4'd8,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd6,4'd4,4'd0};
            8'h07:board={4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd2,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h08:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd2,4'd1,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0};
            8'h09:board={4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0};
            8'h0a:board={4'd1,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd0,4'd5,4'd3,4'd0,4'd0,4'd4,4'd3,4'd0,4'd5,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd5,4'd8,4'd0,4'd7,4'd0,4'd0};
            8'h0b:board={4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd8,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd6,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h0c:board={4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd8,4'd5,4'd0,4'd1,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3};
            8'h0d:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd5,4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0};
            8'h0e:board={4'd0,4'd0,4'd2,4'd0,4'd4,4'd5,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd6,4'd1,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0};
            8'h0f:board={4'd0,4'd0,4'd7,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd2,4'd4,4'd0,4'd6,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0};
            8'h10:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd3,4'd6,4'd1,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0};
            8'h11:board={4'd0,4'd6,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd2,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd7,4'd8};
            8'h12:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd1,4'd0,4'd9,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd5,4'd8,4'd0,4'd0,4'd0};
            8'h13:board={4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd9,4'd7,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0};
            8'h14:board={4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd1};
            8'h15:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0};
            8'h16:board={4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd4,4'd9,4'd0,4'd7,4'd5,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0};
            8'h17:board={4'd0,4'd3,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd1,4'd0,4'd2,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd7,4'd8,4'd0,4'd8,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd4,4'd1,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h18:board={4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd4,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd6,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd4,4'd0,4'd0};
            8'h19:board={4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd9,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3};
            8'h1a:board={4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd2,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd6,4'd2,4'd0,4'd0};
            8'h1b:board={4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd1,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd2,4'd5,4'd0,4'd7,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h1c:board={4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h1d:board={4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd9,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4};
            8'h1e:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd4,4'd3,4'd6,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd4,4'd0};
            8'h1f:board={4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd1,4'd0,4'd7,4'd8,4'd0,4'd2,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd6,4'd8,4'd5,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h20:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd2,4'd5,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd7,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0};
            8'h21:board={4'd8,4'd7,4'd0,4'd0,4'd0,4'd1,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd5,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9};
            8'h22:board={4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd3,4'd5,4'd0,4'd4,4'd6,4'd0,4'd9,4'd4,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3};
            8'h23:board={4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd5,4'd0,4'd6,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd1,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd7,4'd6};
            8'h24:board={4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd8,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h25:board={4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd7,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h26:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0};
            8'h27:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd8,4'd4,4'd3,4'd1,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0};
            8'h28:board={4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd5,4'd0,4'd0,4'd8,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd2,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0};
            8'h29:board={4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9};
            8'h2a:board={4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd1,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7,4'd3,4'd0,4'd0};
            8'h2b:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd9,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd8,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0};
            8'h2c:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd6,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3,4'd8,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd4,4'd9,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0};
            8'h2d:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd8,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5};
            8'h2e:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd8,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd8,4'd4,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd3};
            8'h2f:board={4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd7,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd6,4'd0,4'd1,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0};
            8'h30:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd4,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd9,4'd1,4'd8,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0};
            8'h31:board={4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd4,4'd2,4'd0,4'd9,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd4};
            8'h32:board={4'd4,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd2,4'd9,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4};
            8'h33:board={4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd5,4'd7,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd4,4'd8,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd3,4'd0};
            8'h34:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd5,4'd6,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd6,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0};
            8'h35:board={4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h36:board={4'd0,4'd1,4'd3,4'd4,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3};
            8'h37:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd3,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd7,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd9,4'd4,4'd0};
            8'h38:board={4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd3,4'd0,4'd8,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0};
            8'h39:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd6,4'd3,4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0};
            8'h3a:board={4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd8,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'h3b:board={4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd3,4'd1,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'h3c:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd3,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd1,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd2,4'd0,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h3d:board={4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd7,4'd0,4'd0,4'd4,4'd2,4'd6,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd5,4'd0,4'd4,4'd7,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h3e:board={4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd4,4'd0,4'd2,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd2,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd8,4'd0};
            8'h3f:board={4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0};
            8'h40:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd8,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd6,4'd0,4'd2,4'd0,4'd0,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd1,4'd0,4'd0,4'd4,4'd5,4'd0,4'd6,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0};
            8'h41:board={4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd7,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h42:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd8,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6};
            8'h43:board={4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd5,4'd7,4'd0,4'd4,4'd0,4'd1,4'd1,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd7,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h44:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd3,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd4,4'd0};
            8'h45:board={4'd0,4'd0,4'd1,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd2,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd6,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'h46:board={4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd9,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd8,4'd3,4'd9,4'd0,4'd2,4'd0,4'd4,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd1,4'd8,4'd0,4'd2,4'd6,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd0};
            8'h47:board={4'd6,4'd0,4'd0,4'd2,4'd9,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd1,4'd0,4'd7,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6};
            8'h48:board={4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd6,4'd7,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0};
            8'h49:board={4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd2,4'd4,4'd0,4'd0,4'd0,4'd9,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd7,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd5,4'd8,4'd3,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0};
            8'h4a:board={4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd3,4'd0,4'd1,4'd8,4'd2,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd7,4'd3,4'd0,4'd2,4'd8,4'd0};
            8'h4b:board={4'd0,4'd0,4'd1,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd8,4'd6,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h4c:board={4'd0,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd5,4'd0,4'd2,4'd3,4'd0,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd4,4'd3,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd7};
            8'h4d:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd3,4'd0,4'd6,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h4e:board={4'd0,4'd4,4'd0,4'd5,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd2,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd4,4'd5,4'd4,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0};
            8'h4f:board={4'd5,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd4,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'h50:board={4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd3,4'd1,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd1,4'd7,4'd0,4'd1,4'd0,4'd7,4'd0,4'd5,4'd0,4'd0,4'd8,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd0,4'd3,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd9,4'd0,4'd0};
            8'h51:board={4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0};
            8'h52:board={4'd0,4'd1,4'd8,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd9,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0};
            8'h53:board={4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd6,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd7,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0};
            8'h54:board={4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd2,4'd0,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd7,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6};
            8'h55:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd2,4'd0,4'd4,4'd8,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0};
            8'h56:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd0,4'd0};
            8'h57:board={4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd0,4'd3,4'd7,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd9,4'd8};
            8'h58:board={4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0};
            8'h59:board={4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd9,4'd0,4'd0,4'd4,4'd1,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0};
            8'h5a:board={4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd9,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd5,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0};
            8'h5b:board={4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd6,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd4,4'd9,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h5c:board={4'd1,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd5};
            8'h5d:board={4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd6,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd1,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5};
            8'h5e:board={4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd3,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd9,4'd1,4'd8,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0};
            8'h5f:board={4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd7,4'd2,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd1,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1};
            8'h60:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd6,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd7,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd7,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3};
            8'h61:board={4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd1};
            8'h62:board={4'd7,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd6,4'd4,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0,4'd0};
            8'h63:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd4,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd6,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd7,4'd6,4'd0,4'd2,4'd0,4'd9,4'd8,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3};
            8'h64:board={4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd6,4'd4,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h65:board={4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd6,4'd0,4'd0,4'd7,4'd2,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h66:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd4,4'd0,4'd3,4'd0,4'd1,4'd9,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0};
            8'h67:board={4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd7,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd4,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h68:board={4'd6,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h69:board={4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd4,4'd1,4'd8,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd7,4'd6,4'd8,4'd0,4'd0,4'd4,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6};
            8'h6a:board={4'd0,4'd7,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd9};
            8'h6b:board={4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd8,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd3,4'd6,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h6c:board={4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd2,4'd0,4'd4,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd2,4'd0,4'd6,4'd0,4'd0,4'd7,4'd6,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd8,4'd1};
            8'h6d:board={4'd9,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd2,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd5,4'd7,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1};
            8'h6e:board={4'd6,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd2,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0};
            8'h6f:board={4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd3,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0};
            8'h70:board={4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd4,4'd8,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd2,4'd0,4'd5,4'd7,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0};
            8'h71:board={4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h72:board={4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd7,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0};
            8'h73:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd2,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0};
            8'h74:board={4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd4,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd9,4'd2,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h75:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd5,4'd4,4'd0,4'd2,4'd0,4'd8,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd9,4'd2};
            8'h76:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd8,4'd5,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd9,4'd2,4'd8,4'd0,4'd0,4'd5};
            8'h77:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd8,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd6};
            8'h78:board={4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd3,4'd1,4'd9,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd2,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd6,4'd4,4'd0};
            8'h79:board={4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0};
            8'h7a:board={4'd0,4'd0,4'd0,4'd9,4'd7,4'd3,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd6,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd8,4'd2,4'd5,4'd0,4'd0,4'd3,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9};
            8'h7b:board={4'd1,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd0,4'd8,4'd6,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd5,4'd9,4'd0,4'd7,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h7c:board={4'd2,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0};
            8'h7d:board={4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd8,4'd0,4'd9,4'd7,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd1,4'd0,4'd0,4'd0};
            8'h7e:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd0,4'd2,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd0,4'd8,4'd0,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd1,4'd9,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h7f:board={4'd0,4'd6,4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd4,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd5};
            8'h80:board={4'd7,4'd0,4'd3,4'd0,4'd0,4'd8,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd9,4'd3,4'd8,4'd0};
            8'h81:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd6,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd2,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd5,4'd6,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h82:board={4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd3,4'd0,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd4,4'd4,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h83:board={4'd7,4'd3,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd5,4'd0,4'd4,4'd6,4'd0};
            8'h84:board={4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd9,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd3};
            8'h85:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd4,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0};
            8'h86:board={4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd7,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h87:board={4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd9,4'd6,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd6,4'd0};
            8'h88:board={4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd7,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd5,4'd6,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0};
            8'h89:board={4'd5,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd1,4'd8,4'd2,4'd3,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd5,4'd0,4'd1,4'd8,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h8a:board={4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd1,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd1,4'd0,4'd0,4'd0,4'd8,4'd3,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'h8b:board={4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd1,4'd6,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd4,4'd0,4'd9,4'd6,4'd0,4'd0};
            8'h8c:board={4'd2,4'd6,4'd0,4'd0,4'd0,4'd9,4'd1,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0};
            8'h8d:board={4'd2,4'd1,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd5,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd0,4'd5,4'd8,4'd0,4'd7,4'd6,4'd0,4'd0,4'd4};
            8'h8e:board={4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd9,4'd2,4'd0,4'd0,4'd0,4'd0};
            8'h8f:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd1,4'd6,4'd4,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd2,4'd0};
            8'h90:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd2,4'd5,4'd8,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0};
            8'h91:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd5,4'd3,4'd8,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd3,4'd4,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd0,4'd5,4'd7,4'd0};
            8'h92:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd4,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd3,4'd8,4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0};
            8'h93:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd6,4'd3,4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0};
            8'h94:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd1,4'd4,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd2,4'd3,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd2,4'd7,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0};
            8'h95:board={4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd5,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd9,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd6,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0};
            8'h96:board={4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd4,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0};
            8'h97:board={4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd1,4'd0,4'd0,4'd2,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd7,4'd5,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd4,4'd5,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0};
            8'h98:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd4,4'd0,4'd3,4'd6,4'd5,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd2,4'd0,4'd9,4'd0,4'd0};
            8'h99:board={4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd8,4'd7,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0};
            8'h9a:board={4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0};
            8'h9b:board={4'd4,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0};
            8'h9c:board={4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd6,4'd1,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd3,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0};
            8'h9d:board={4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd3,4'd0,4'd8,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0};
            8'h9e:board={4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd5,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            8'h9f:board={4'd0,4'd0,4'd6,4'd0,4'd4,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd2,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd1,4'd9,4'd3,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd7,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'ha0:board={4'd2,4'd9,4'd0,4'd6,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd5,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'ha1:board={4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd7,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd3,4'd0,4'd0};
            8'ha2:board={4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd0,4'd0,4'd8};
            8'ha3:board={4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd8,4'd5,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd5,4'd2,4'd0,4'd9,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd8,4'd1,4'd0,4'd6,4'd0,4'd0,4'd1,4'd6,4'd9,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'ha4:board={4'd2,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd4,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd8,4'd9,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'ha5:board={4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd8,4'd8,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd8,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd0};
            8'ha6:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd4,4'd0,4'd0,4'd4,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd8,4'd0,4'd9,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0};
            8'ha7:board={4'd1,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0};
            8'ha8:board={4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd4,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd7,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'ha9:board={4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd8,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd4,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd3,4'd4,4'd0,4'd0,4'd0,4'd6};
            8'haa:board={4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd2,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd9,4'd0,4'd1,4'd0,4'd3,4'd2,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0};
            8'hab:board={4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd3,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd9,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8};
            8'hac:board={4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd8,4'd0,4'd2,4'd9,4'd0,4'd0};
            8'had:board={4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd2,4'd0,4'd3,4'd8,4'd0,4'd6,4'd0,4'd5,4'd6,4'd0,4'd9,4'd5,4'd1,4'd0,4'd7,4'd0,4'd0};
            8'hae:board={4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd3,4'd0,4'd8,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd8,4'd6,4'd4,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd9,4'd7};
            8'haf:board={4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd2,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd7,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd2,4'd7,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0};
            8'hb0:board={4'd0,4'd4,4'd0,4'd2,4'd9,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd8,4'd6,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd9,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd9,4'd0,4'd0};
            8'hb1:board={4'd0,4'd7,4'd0,4'd0,4'd2,4'd1,4'd5,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd3};
            8'hb2:board={4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd2,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd3,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd3,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hb3:board={4'd7,4'd0,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd8,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0};
            8'hb4:board={4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd5};
            8'hb5:board={4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd9,4'd0,4'd2,4'd5,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7};
            8'hb6:board={4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd1,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0};
            8'hb7:board={4'd0,4'd0,4'd7,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd2,4'd4,4'd0,4'd6,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0};
            8'hb8:board={4'd2,4'd0,4'd0,4'd0,4'd6,4'd4,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd7,4'd9,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0};
            8'hb9:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd0,4'd1,4'd9,4'd7,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd2,4'd4,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0};
            8'hba:board={4'd4,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd7,4'd3,4'd0,4'd0,4'd4,4'd0,4'd7,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd7,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd6,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0};
            8'hbb:board={4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd3,4'd0,4'd4,4'd8,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd6,4'd0};
            8'hbc:board={4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0};
            8'hbd:board={4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd9,4'd4,4'd0,4'd2,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0};
            8'hbe:board={4'd0,4'd0,4'd0,4'd5,4'd4,4'd8,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd9,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7};
            8'hbf:board={4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd3,4'd5,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd7,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hc0:board={4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0};
            8'hc1:board={4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd1,4'd0,4'd6,4'd0,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0};
            8'hc2:board={4'd0,4'd0,4'd0,4'd4,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd7,4'd1,4'd0,4'd9,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hc3:board={4'd4,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd9,4'd0,4'd9,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd8,4'd0,4'd7,4'd8,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hc4:board={4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd7,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0};
            8'hc5:board={4'd5,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd7,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd4,4'd2,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0};
            8'hc6:board={4'd3,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd2,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd4,4'd0,4'd1,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1};
            8'hc7:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0};
            8'hc8:board={4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd1,4'd6,4'd0,4'd2,4'd0,4'd5,4'd1,4'd0,4'd0,4'd4,4'd9,4'd0,4'd3,4'd0,4'd8,4'd2,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd1};
            8'hc9:board={4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd3,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd4,4'd0,4'd0,4'd3,4'd0,4'd1,4'd2};
            8'hca:board={4'd0,4'd3,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5};
            8'hcb:board={4'd0,4'd0,4'd1,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd5,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0};
            8'hcc:board={4'd0,4'd7,4'd8,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd9,4'd0,4'd4,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd8,4'd4,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0};
            8'hcd:board={4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd5,4'd3,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd7,4'd7,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0};
            8'hce:board={4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd7,4'd0,4'd0,4'd1,4'd8,4'd2,4'd4,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0};
            8'hcf:board={4'd3,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd2,4'd6,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd1,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd8};
            8'hd0:board={4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd4,4'd8,4'd0,4'd2,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd5,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd2,4'd0,4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0};
            8'hd1:board={4'd9,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd7,4'd9,4'd0,4'd5,4'd0,4'd0,4'd5,4'd8,4'd9,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0};
            8'hd2:board={4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd2,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd8,4'd0,4'd0};
            8'hd3:board={4'd0,4'd4,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd1,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd8,4'd0,4'd0,4'd9,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hd4:board={4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd8,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0};
            8'hd5:board={4'd0,4'd9,4'd1,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd8,4'd6,4'd3,4'd2,4'd0,4'd0,4'd0,4'd7,4'd3,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd2,4'd3,4'd0};
            8'hd6:board={4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd1,4'd0,4'd1,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd5,4'd4,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd5,4'd0,4'd8,4'd0,4'd6,4'd0,4'd4,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hd7:board={4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd5,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd1,4'd0,4'd8,4'd7,4'd0,4'd5,4'd8,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hd8:board={4'd7,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd7,4'd4,4'd7,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hd9:board={4'd2,4'd8,4'd9,4'd3,4'd0,4'd1,4'd0,4'd7,4'd0,4'd7,4'd4,4'd0,4'd0,4'd2,4'd0,4'd5,4'd1,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd2,4'd0,4'd5,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd8,4'd7,4'd0,4'd0,4'd4,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hda:board={4'd3,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd9,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2};
            8'hdb:board={4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd2,4'd0,4'd2,4'd5,4'd4,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd4,4'd1,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0};
            8'hdc:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd6,4'd4,4'd0,4'd0,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd3,4'd7,4'd5,4'd0,4'd0,4'd1,4'd8,4'd7,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hdd:board={4'd4,4'd0,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd4,4'd2,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hde:board={4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd5,4'd0,4'd0,4'd7,4'd1,4'd5,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hdf:board={4'd0,4'd8,4'd7,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd4,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd4,4'd0,4'd8,4'd0,4'd0};
            8'he0:board={4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd3,4'd8,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd6,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd0,4'd8,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0};
            8'he1:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd5,4'd1,4'd8,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd6,4'd0,4'd6,4'd0,4'd8,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd0,4'd2,4'd0,4'd0};
            8'he2:board={4'd0,4'd7,4'd0,4'd0,4'd1,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd8,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0};
            8'he3:board={4'd0,4'd2,4'd8,4'd0,4'd3,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd4,4'd0,4'd2};
            8'he4:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd5,4'd9,4'd0};
            8'he5:board={4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd2,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd5,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6};
            8'he6:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd1,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd2,4'd7};
            8'he7:board={4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd7,4'd2};
            8'he8:board={4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd7,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'he9:board={4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd1,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd5,4'd8,4'd4};
            8'hea:board={4'd0,4'd0,4'd3,4'd4,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd2,4'd5,4'd0,4'd6,4'd0,4'd9,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd8,4'd2,4'd0,4'd4,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'heb:board={4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd0,4'd3,4'd8,4'd7,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0};
            8'hec:board={4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd8,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd7,4'd0};
            8'hed:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd5,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd4,4'd0,4'd5,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd2,4'd0,4'd6,4'd4,4'd0,4'd0,4'd0};
            8'hee:board={4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd9,4'd0,4'd0,4'd5,4'd3,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd2};
            8'hef:board={4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd7,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hf0:board={4'd0,4'd4,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0};
            8'hf1:board={4'd0,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0};
            8'hf2:board={4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd2,4'd5,4'd5,4'd3,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd4,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0};
            8'hf3:board={4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd6,4'd7,4'd4,4'd0,4'd7,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd4,4'd8,4'd2,4'd0,4'd7,4'd0,4'd0};
            8'hf4:board={4'd0,4'd9,4'd0,4'd3,4'd2,4'd0,4'd0,4'd0,4'd6,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0};
            8'hf5:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd3,4'd9,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd1,4'd5,4'd0,4'd4,4'd0,4'd6,4'd2,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd9,4'd0,4'd4,4'd0,4'd0,4'd8,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hf6:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd1,4'd4,4'd0,4'd3,4'd2,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd8,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0};
            8'hf7:board={4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd9,4'd6,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd7,4'd4,4'd3,4'd8,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0};
            8'hf8:board={4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd5,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            8'hf9:board={4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd7,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd3,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd2,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0};
            8'hfa:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd2,4'd5,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd5,4'd2,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0};
            8'hfb:board={4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd5,4'd0,4'd8,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd9,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd4,4'd7,4'd0,4'd3};
            8'hfc:board={4'd7,4'd5,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd9,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd8,4'd0,4'd2,4'd0,4'd9,4'd0,4'd0};
            8'hfd:board={4'd7,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd1,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd1,4'd0,4'd8,4'd2,4'd0,4'd0};
            8'hfe:board={4'd3,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd5,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd8,4'd0,4'd6,4'd0,4'd3,4'd4,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4};
        endcase
    end
endmodule