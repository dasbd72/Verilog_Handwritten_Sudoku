`timescale 1ps/1ps
module SudokuGenerator #(
    parameter size = 4'd9,
    parameter bit = 4'd4
    ) (
    input [15:0] random,
    output reg [81*4-1:0] board,
    output wire [81-1:0]  board_blank
    );
    
    genvar i;
    generate
        for(i = 0; i < 81; i = i + 1) begin
            assign board_blank[i] = board[(i+1)*bit-1-:bit] == 4'd0;
        end
    endgenerate

    always @(*) begin
        case (random[5:0])
            6'h00:board={4'd8,4'd0,4'd4,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd4,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd7,4'd7,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0};
            6'h01:board={4'd3,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd4,4'd9,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2};
            6'h02:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd2,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd9,4'd2,4'd3,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd4,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0};
            6'h03:board={4'd2,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd4,4'd0,4'd9,4'd0,4'd5,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd3,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0};
            6'h04:board={4'd0,4'd9,4'd0,4'd2,4'd0,4'd4,4'd5,4'd0,4'd0,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd9,4'd5,4'd0,4'd0,4'd8,4'd0,4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd9};
            6'h05:board={4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd6,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h06:board={4'd6,4'd1,4'd0,4'd8,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd6,4'd4,4'd0};
            6'h07:board={4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd2,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h08:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd8,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd2,4'd1,4'd0,4'd9,4'd3,4'd0,4'd0,4'd0};
            6'h09:board={4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0};
            6'h0a:board={4'd1,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd0,4'd5,4'd3,4'd0,4'd0,4'd4,4'd3,4'd0,4'd5,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd5,4'd8,4'd0,4'd7,4'd0,4'd0};
            6'h0b:board={4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd8,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd0,4'd6,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h0c:board={4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd8,4'd5,4'd0,4'd1,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3};
            6'h0d:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd5,4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd1,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0};
            6'h0e:board={4'd0,4'd0,4'd2,4'd0,4'd4,4'd5,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd6,4'd1,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd4,4'd0};
            6'h0f:board={4'd0,4'd0,4'd7,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd2,4'd4,4'd0,4'd6,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0};
            6'h10:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd3,4'd0,4'd2,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd3,4'd6,4'd1,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0};
            6'h11:board={4'd0,4'd6,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd2,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd7,4'd8};
            6'h12:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd1,4'd0,4'd9,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd5,4'd8,4'd0,4'd0,4'd0};
            6'h13:board={4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd3,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd9,4'd7,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd2,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0};
            6'h14:board={4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd3,4'd0,4'd4,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd1};
            6'h15:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd1,4'd0,4'd0};
            6'h16:board={4'd0,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd3,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd0,4'd4,4'd9,4'd0,4'd7,4'd5,4'd3,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd8,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0};
            6'h17:board={4'd0,4'd3,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd3,4'd1,4'd0,4'd2,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd7,4'd8,4'd0,4'd8,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd8,4'd0,4'd0,4'd4,4'd1,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h18:board={4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd4,4'd3,4'd0,4'd7,4'd0,4'd0,4'd0,4'd6,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd6,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd8,4'd4,4'd0,4'd0};
            6'h19:board={4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd9,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3};
            6'h1a:board={4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd2,4'd4,4'd0,4'd0,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd2,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd0,4'd6,4'd2,4'd0,4'd0};
            6'h1b:board={4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd1,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd2,4'd5,4'd0,4'd7,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd9,4'd0,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd6,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h1c:board={4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd9,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            6'h1d:board={4'd0,4'd6,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd9,4'd5,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4};
            6'h1e:board={4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd4,4'd3,4'd6,4'd0,4'd1,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd3,4'd0,4'd0,4'd2,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd3,4'd0,4'd4,4'd0};
            6'h1f:board={4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd9,4'd1,4'd0,4'd7,4'd8,4'd0,4'd2,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd6,4'd8,4'd5,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h20:board={4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd2,4'd5,4'd9,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd0,4'd0,4'd8,4'd7,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0};
            6'h21:board={4'd8,4'd7,4'd0,4'd0,4'd0,4'd1,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd5,4'd0,4'd8,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9};
            6'h22:board={4'd1,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd0,4'd0,4'd0,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd3,4'd5,4'd0,4'd4,4'd6,4'd0,4'd9,4'd4,4'd6,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3};
            6'h23:board={4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd4,4'd5,4'd0,4'd6,4'd0,4'd0,4'd3,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd1,4'd1,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd7,4'd6};
            6'h24:board={4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd7,4'd0,4'd9,4'd0,4'd4,4'd0,4'd0,4'd8,4'd6,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd2,4'd5,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd1,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2};
            6'h25:board={4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd0,4'd7,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd7,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h26:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd6,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd2,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd6,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0};
            6'h27:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd7,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd7,4'd0,4'd8,4'd4,4'd3,4'd1,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0};
            6'h28:board={4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd7,4'd5,4'd0,4'd0,4'd8,4'd9,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd7,4'd2,4'd0,4'd1,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd2,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd6,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd1,4'd0};
            6'h29:board={4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd4,4'd1,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd9,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd9};
            6'h2a:board={4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd9,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd2,4'd1,4'd9,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd7,4'd3,4'd0,4'd0};
            6'h2b:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd6,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd9,4'd2,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd8,4'd9,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0};
            6'h2c:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd6,4'd9,4'd0,4'd0,4'd2,4'd0,4'd0,4'd3,4'd8,4'd0,4'd2,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd6,4'd1,4'd0,4'd4,4'd9,4'd0,4'd0,4'd3,4'd0,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0};
            6'h2d:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd4,4'd9,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd8,4'd0,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd2,4'd0,4'd0,4'd8,4'd2,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5};
            6'h2e:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd8,4'd1,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd8,4'd4,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd3};
            6'h2f:board={4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd7,4'd0,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd6,4'd0,4'd1,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd8,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0};
            6'h30:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd9,4'd0,4'd4,4'd2,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd3,4'd4,4'd0,4'd0,4'd8,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd9,4'd1,4'd8,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd9,4'd4,4'd0};
            6'h31:board={4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd6,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd6,4'd4,4'd2,4'd0,4'd9,4'd3,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd0,4'd8,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd4};
            6'h32:board={4'd4,4'd6,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd3,4'd0,4'd5,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd3,4'd0,4'd0,4'd0,4'd2,4'd9,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd8,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd2,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd4};
            6'h33:board={4'd0,4'd0,4'd1,4'd0,4'd9,4'd0,4'd5,4'd7,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd3,4'd0,4'd0,4'd0,4'd9,4'd7,4'd0,4'd0,4'd4,4'd8,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd5,4'd8,4'd0,4'd0,4'd0,4'd3,4'd0};
            6'h34:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd2,4'd5,4'd6,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd3,4'd2,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd0,4'd9,4'd6,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd4,4'd0,4'd0,4'd6,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0};
            6'h35:board={4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd4,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd3,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd1,4'd0,4'd0,4'd0,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd7,4'd1,4'd0,4'd0,4'd0,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h36:board={4'd0,4'd1,4'd3,4'd4,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd2,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd3,4'd1,4'd0,4'd0,4'd0,4'd0,4'd9,4'd1,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd3};
            6'h37:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd2,4'd3,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd7,4'd1,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd8,4'd3,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd9,4'd4,4'd0};
            6'h38:board={4'd0,4'd0,4'd0,4'd7,4'd8,4'd0,4'd0,4'd3,4'd0,4'd8,4'd1,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd6,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd1,4'd0,4'd0,4'd6,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd0,4'd5,4'd0};
            6'h39:board={4'd6,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd2,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd3,4'd6,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd0,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd5,4'd7,4'd0,4'd0,4'd6,4'd3,4'd7,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd3,4'd0,4'd1,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0};
            6'h3a:board={4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd0,4'd9,4'd0,4'd1,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd8,4'd6,4'd0,4'd3,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd5,4'd0,4'd7,4'd0,4'd8,4'd6,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8};
            6'h3b:board={4'd0,4'd8,4'd0,4'd3,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd2,4'd0,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd8,4'd0,4'd0,4'd0,4'd0,4'd1,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd9,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd2,4'd3,4'd1,4'd6,4'd4,4'd0,4'd0,4'd0,4'd0,4'd8};
            6'h3c:board={4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd9,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd2,4'd0,4'd0,4'd3,4'd1,4'd7,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd7,4'd0,4'd0,4'd0,4'd0,4'd9,4'd2,4'd1,4'd5,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd2,4'd0,4'd0,4'd8,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h3d:board={4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd8,4'd7,4'd0,4'd0,4'd4,4'd2,4'd6,4'd0,4'd0,4'd0,4'd3,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd5,4'd0,4'd4,4'd7,4'd0,4'd0,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd1,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd9,4'd0,4'd0,4'd7,4'd0,4'd2,4'd0,4'd5,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0};
            6'h3e:board={4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd0,4'd8,4'd4,4'd0,4'd2,4'd0,4'd5,4'd7,4'd0,4'd0,4'd0,4'd3,4'd0,4'd7,4'd0,4'd2,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd4,4'd2,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd5,4'd1,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd9,4'd2,4'd0,4'd1,4'd0,4'd7,4'd0,4'd0,4'd4,4'd0,4'd8,4'd0};
            6'h3f:board={4'd1,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd4,4'd0,4'd6,4'd0,4'd0,4'd8,4'd0,4'd0,4'd3,4'd0,4'd0,4'd7,4'd0,4'd4,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd3,4'd0,4'd6,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd9,4'd0,4'd2,4'd0,4'd0,4'd0,4'd6,4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd2,4'd0,4'd0,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd0};
        endcase
    end
endmodule