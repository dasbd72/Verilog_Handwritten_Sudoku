/*
    clk : posedge clock signal
    rst : posedge reset signal
    start : req 1 cycle signal
    layer_input : req 64 cycle
    layer_0 : last until next start signal
    finish : last 1 cycle
 */
module Dense_0(
    input  wire clk, 
    input  wire rst,
    input  wire start,
    input  wire [28*28 - 1:0] layer_input,
    output reg  [16*64 - 1:0] layer_0,
    output reg  finish
    );
    localparam HEIGHT = 784;
    localparam WIDTH = 64;
    localparam [802815:0] kernel_0 = {16'h0069,16'h00a5,-16'h005d,-16'h0132,16'h004b,-16'h0002,-16'h0077,16'h00da,16'h015c,-16'h0082,-16'h0030,16'h0083,16'h004c,16'h0167,-16'h0056,-16'h0170,-16'h00af,16'h00f8,-16'h0030,16'h0070,-16'h00b2,16'h0185,-16'h0010,16'h0027,-16'h0013,16'h000c,-16'h00a6,-16'h0016,-16'h0035,-16'h0006,-16'h0107,-16'h0096,-16'h0049,-16'h0138,-16'h00f3,-16'h00b7,-16'h011e,-16'h00a9,16'h01b8,-16'h00ea,-16'h0089,16'h014a,-16'h0006,16'h01f8,16'h008e,16'h00bb,-16'h00d8,-16'h00a7,16'h01f3,16'h003f,16'h00e5,-16'h0098,-16'h006a,-16'h0053,-16'h0170,16'h005e,16'h0162,-16'h01db,16'h0094,16'h0062,16'h0190,16'h0038,-16'h0068,-16'h0121,-16'h0058,16'h0044,-16'h006e,-16'h00d9,16'h010b,16'h0050,16'h003f,16'h0067,16'h002b,-16'h0174,-16'h0009,-16'h0012,16'h0015,16'h0187,-16'h0043,-16'h01ee,-16'h003c,16'h00ac,-16'h00b1,16'h002e,-16'h0024,16'h00b9,16'h0072,-16'h0044,16'h00a0,16'h008b,-16'h0128,16'h0029,16'h0058,16'h006c,-16'h00b7,-16'h0029,-16'h0025,-16'h0078,-16'h00c4,-16'h0082,-16'h00db,-16'h0026,16'h023b,16'h0030,-16'h0106,16'h014d,-16'h0035,16'h015f,16'h002b,16'h00df,-16'h00cd,-16'h0088,16'h020e,16'h002f,16'h00a1,-16'h008c,-16'h00a2,-16'h0018,-16'h0062,16'h00b7,16'h0116,-16'h020e,16'h008c,16'h002f,16'h0108,-16'h0008,-16'h00d2,-16'h00fe,-16'h00ca,16'h002e,-16'h011a,-16'h00bd,16'h00b5,16'h00e1,16'h000a,-16'h0027,16'h0050,-16'h01f0,16'h0057,16'h004b,-16'h0039,16'h01a4,-16'h000a,-16'h01ed,-16'h0012,16'h011a,-16'h0117,16'h0085,-16'h0081,16'h0062,-16'h0043,-16'h0055,16'h00f2,16'h000a,-16'h0145,16'h002b,16'h004f,16'h000e,-16'h0051,-16'h004b,16'h0040,-16'h00bf,-16'h004b,-16'h0046,-16'h0153,16'h0058,16'h0288,16'h0096,-16'h010c,16'h011b,-16'h0075,16'h01b8,16'h00b5,16'h00e9,-16'h006c,-16'h0038,16'h019b,16'h002d,16'h0118,-16'h00aa,-16'h00b3,-16'h002b,-16'h0085,16'h0026,16'h017a,-16'h0139,16'h00b7,16'h004c,16'h0053,16'h0041,-16'h0169,-16'h015e,-16'h00ba,16'h0063,-16'h01bd,-16'h0072,16'h00b0,16'h012a,16'h0000,16'h000f,16'h000c,-16'h01ad,16'h005a,-16'h0028,-16'h0092,16'h01c1,16'h002f,-16'h0140,16'h0052,16'h0112,-16'h0179,16'h0042,-16'h0002,16'h012c,16'h0048,-16'h0100,16'h011c,16'h0098,-16'h00f9,16'h0031,16'h0036,16'h003f,-16'h003f,-16'h002f,16'h00ee,-16'h0074,-16'h0031,16'h0006,-16'h01dd,-16'h0002,16'h034e,16'h0054,-16'h019a,16'h00ff,16'h0005,16'h01d7,16'h00ee,16'h01a0,-16'h00ec,-16'h0020,16'h01a2,-16'h0064,16'h0111,-16'h00f5,-16'h0197,-16'h0039,-16'h00cd,-16'h0007,16'h00f6,-16'h0028,16'h0084,16'h002b,-16'h0077,16'h004f,-16'h00f5,-16'h01c9,-16'h013f,16'h00ca,-16'h01e7,-16'h0003,16'h01ac,16'h0080,16'h0016,-16'h0043,-16'h0059,-16'h0139,16'h0010,-16'h00ad,-16'h0163,16'h014e,-16'h0021,16'h0000,16'h00be,16'h0025,-16'h01ad,16'h000b,16'h0003,16'h010d,16'h0047,-16'h01ab,16'h00e9,16'h00a8,-16'h009e,16'h0075,16'h007d,16'h0013,-16'h006d,16'h0031,16'h00a4,-16'h004c,-16'h00a0,16'h009d,-16'h0228,16'h0065,16'h0348,16'h002d,-16'h017d,16'h0139,16'h001d,16'h0177,16'h004e,16'h01f0,-16'h00fe,16'h0056,16'h01a9,-16'h0072,16'h00d1,-16'h0170,-16'h01ee,-16'h00a0,-16'h002d,16'h0084,16'h015f,16'h003e,16'h0058,16'h0067,-16'h00ed,-16'h0041,-16'h0081,-16'h01d7,-16'h007c,16'h0126,-16'h027f,-16'h0039,16'h0199,16'h0006,16'h0006,16'h0002,-16'h002c,-16'h0086,16'h004f,-16'h00d8,-16'h01cf,16'h018a,16'h0011,16'h002a,16'h0062,-16'h008c,-16'h01a2,16'h002b,16'h0030,16'h00d7,16'h00b8,-16'h0193,16'h00d8,16'h0060,-16'h0021,16'h007c,16'h003e,16'h0000,-16'h00b5,-16'h0020,16'h008e,-16'h0015,-16'h0140,16'h008b,-16'h01a5,16'h00ae,16'h02c9,-16'h00a2,-16'h01c8,16'h00d6,16'h0051,16'h00b5,16'h0089,16'h0144,-16'h00e9,16'h001b,16'h0087,-16'h00c8,16'h00ac,-16'h012b,-16'h01ee,-16'h0082,-16'h0063,16'h006b,16'h0186,16'h0129,16'h007c,16'h00a9,-16'h009b,-16'h009e,-16'h0085,-16'h0193,16'h0058,16'h0162,-16'h0330,-16'h003e,16'h0237,16'h0016,-16'h001c,16'h002d,-16'h0114,-16'h007b,16'h003d,-16'h0145,-16'h026b,16'h0175,-16'h0023,16'h0067,16'h001b,-16'h013e,-16'h01e0,16'h0049,16'h0080,16'h004e,16'h00bc,-16'h0202,-16'h007e,16'h0063,16'h003f,16'h0068,16'h002a,-16'h005a,-16'h003d,16'h0020,16'h0070,16'h009f,-16'h012d,16'h00a6,-16'h010c,16'h007e,16'h02ed,-16'h0062,-16'h01c1,16'h013e,16'h00a4,16'h00dc,16'h0046,16'h00e1,-16'h017a,16'h0034,-16'h0012,-16'h0105,16'h0066,-16'h01f4,-16'h0119,-16'h00a0,16'h0034,16'h0045,16'h0117,16'h010f,16'h0017,16'h00b6,-16'h0082,-16'h0095,-16'h00d1,-16'h01c7,16'h0035,16'h016a,-16'h041e,-16'h0071,16'h0268,16'h002f,-16'h0028,16'h0098,-16'h00dc,-16'h0077,-16'h000d,-16'h0144,-16'h01d7,16'h00cb,16'h004f,16'h0083,-16'h0020,-16'h00fe,-16'h014d,16'h0083,16'h00a6,16'h008b,16'h00d8,-16'h019d,-16'h0224,16'h00c3,16'h000e,16'h00f0,16'h0065,-16'h0036,16'h001a,-16'h0083,16'h00f4,16'h006e,-16'h013d,16'h00b6,-16'h009f,16'h0081,16'h027a,-16'h006c,-16'h02e3,16'h01b4,16'h0129,-16'h000f,16'h0081,16'h006f,-16'h0150,-16'h004b,16'h007e,-16'h01e8,-16'h0037,-16'h0249,16'h0026,-16'h0030,16'h0081,16'h00d2,16'h0089,16'h010b,16'h0089,16'h00a7,16'h0030,-16'h0050,-16'h0089,-16'h016a,16'h0041,16'h01ae,-16'h0436,16'h0032,16'h0236,16'h0082,-16'h0043,16'h003f,-16'h00a7,-16'h004c,16'h0003,-16'h013f,-16'h0190,16'h0075,16'h0040,16'h0011,16'h0027,-16'h012d,-16'h0111,16'h00aa,16'h007f,16'h00a8,16'h0163,-16'h01d0,-16'h0359,16'h0121,-16'h0033,16'h007b,16'h011c,-16'h006c,16'h00dd,-16'h00aa,16'h0175,16'h004b,-16'h01b0,16'h0082,16'h001a,-16'h0083,16'h024f,-16'h0078,-16'h029e,16'h016e,16'h0088,16'h0001,16'h0078,16'h0058,-16'h01bf,-16'h007b,-16'h003c,-16'h0282,16'h001c,-16'h01f7,-16'h0057,-16'h0044,16'h000d,16'h0035,16'h0033,16'h017a,16'h001f,16'h0105,16'h005d,-16'h007b,-16'h0055,-16'h014a,-16'h000e,16'h0107,-16'h0371,16'h0039,16'h020b,16'h0083,-16'h0040,-16'h0054,-16'h0098,-16'h001f,-16'h0098,-16'h00e8,-16'h00b6,-16'h0007,-16'h0052,-16'h0012,-16'h0007,-16'h0118,-16'h00e6,16'h0011,16'h0051,-16'h0017,16'h01a4,-16'h0195,-16'h03e2,16'h0128,-16'h00ae,16'h0033,16'h0128,-16'h0062,16'h005b,-16'h0068,16'h01db,16'h0049,-16'h0136,-16'h008c,16'h007f,-16'h00c1,16'h025c,-16'h0060,-16'h0334,16'h0132,16'h003c,16'h0023,16'h0079,16'h0060,-16'h0246,-16'h00e5,16'h001c,-16'h01de,16'h0016,-16'h0136,16'h004d,-16'h0029,16'h007b,16'h00e5,16'h0120,16'h01a4,-16'h0041,16'h00c4,16'h0080,-16'h004d,16'h0071,-16'h00e9,16'h0074,16'h00c7,-16'h033f,-16'h0030,16'h0211,16'h000b,-16'h00ff,-16'h0056,-16'h000e,16'h0059,16'h0049,-16'h00fc,16'h003d,-16'h00ab,16'h0038,-16'h00b3,16'h00f5,-16'h0184,-16'h004d,16'h008e,16'h007a,-16'h0015,16'h013d,-16'h017d,-16'h044e,16'h00f8,16'h0002,16'h00c4,16'h00ee,-16'h00a6,16'h0047,-16'h00f6,16'h01ad,16'h0010,-16'h01bf,16'h0000,16'h00cf,-16'h0098,16'h0228,-16'h0005,-16'h03a1,16'h0175,-16'h000e,16'h0069,16'h00b5,-16'h001c,-16'h0306,-16'h01cb,16'h0013,-16'h0186,-16'h0036,-16'h00d2,-16'h0037,16'h0071,16'h00ba,16'h00de,16'h0046,16'h0193,-16'h0089,16'h0150,16'h0057,-16'h0104,-16'h001d,-16'h00c2,-16'h002d,16'h006f,-16'h029f,-16'h0061,16'h022a,16'h0000,-16'h0105,-16'h0025,-16'h0020,16'h018c,-16'h0014,-16'h0082,16'h00c8,-16'h010a,16'h0053,-16'h0173,16'h0092,-16'h0107,-16'h006b,16'h001e,-16'h0024,16'h0009,16'h00e5,-16'h01aa,-16'h042c,16'h00be,-16'h000f,16'h0063,16'h013f,-16'h009b,-16'h0044,-16'h003e,16'h016b,16'h002b,-16'h01cf,-16'h008e,16'h0132,-16'h00ad,16'h01ac,16'h0063,-16'h0391,16'h0150,16'h002c,-16'h0002,16'h001d,-16'h00c7,-16'h0386,-16'h02bf,16'h0068,-16'h024f,-16'h0043,-16'h0001,-16'h0007,16'h004e,16'h005c,16'h006f,16'h000d,16'h0063,-16'h00b3,16'h0127,-16'h002d,-16'h004b,16'h000b,-16'h00e7,16'h001f,16'h00fd,-16'h0281,-16'h0165,16'h01cb,-16'h0021,-16'h016e,16'h005e,16'h0043,16'h01f6,16'h0083,-16'h001e,16'h00bc,-16'h0094,-16'h0005,-16'h0157,16'h00ef,-16'h0121,-16'h00a4,16'h0000,-16'h0011,16'h0052,16'h004f,-16'h01bd,-16'h03ae,16'h00c4,-16'h0004,16'h0076,16'h00b9,-16'h008b,-16'h0083,-16'h00dc,16'h018c,16'h004b,-16'h014c,-16'h0040,16'h0172,-16'h000b,16'h020d,16'h0067,-16'h02af,16'h01bc,16'h0059,16'h0045,16'h009c,-16'h00b4,-16'h0438,-16'h0343,16'h0046,-16'h0217,-16'h0085,-16'h008c,-16'h003b,16'h00c9,-16'h0018,16'h0088,-16'h0047,-16'h011c,-16'h00ad,16'h016a,-16'h004e,-16'h005c,16'h003a,-16'h009b,-16'h0002,16'h00bd,-16'h01be,-16'h0284,16'h01d6,-16'h0053,-16'h0112,16'h0050,16'h002e,16'h023d,16'h008d,-16'h0023,16'h0101,-16'h0109,16'h0075,-16'h005b,16'h00dd,-16'h0100,-16'h0030,16'h009e,-16'h0019,16'h0053,16'h0027,-16'h01dc,-16'h028e,16'h011b,-16'h000c,16'h00f9,16'h0072,-16'h0094,-16'h00c0,16'h0011,16'h011a,16'h001e,-16'h00b5,-16'h0087,16'h01ab,16'h002d,16'h01b0,16'h00cf,-16'h0370,16'h017c,16'h00e6,16'h0076,16'h0018,-16'h00f2,-16'h0468,-16'h0406,16'h004d,-16'h025d,-16'h0112,-16'h0030,-16'h00e3,16'h009e,16'h0064,16'h007d,-16'h0074,-16'h0103,-16'h007f,16'h01a0,-16'h00bd,-16'h008d,16'h0045,-16'h00dc,16'h007a,16'h009e,-16'h0114,-16'h0324,16'h0189,-16'h007c,-16'h00e2,16'h0059,-16'h004c,16'h0218,16'h00ad,-16'h0064,16'h0181,-16'h0064,16'h007c,16'h003b,16'h0102,-16'h004e,-16'h003d,-16'h0034,16'h0023,16'h0017,16'h0058,-16'h0165,-16'h0236,16'h00ba,16'h005a,16'h007e,16'h0066,-16'h010f,-16'h0170,16'h0046,16'h0130,-16'h002e,-16'h0051,-16'h004c,16'h0166,16'h005a,16'h01c0,16'h0099,-16'h033b,16'h012c,16'h004f,16'h00bf,16'h00a5,-16'h019a,-16'h04cb,-16'h02fd,16'h0027,-16'h02ec,-16'h00f4,-16'h005a,-16'h0079,16'h0101,16'h00ea,16'h0032,-16'h00b8,-16'h0111,16'h000e,16'h0113,-16'h0030,-16'h00d1,16'h0067,-16'h016c,-16'h0038,16'h00e1,-16'h0137,-16'h02fb,16'h0186,-16'h005c,-16'h00ef,16'h0061,16'h001f,16'h025c,16'h00f7,-16'h0012,16'h0142,16'h001d,16'h00a7,16'h0138,16'h00e7,16'h003b,-16'h00d3,-16'h0044,16'h0001,-16'h0002,-16'h0053,-16'h0109,-16'h016d,-16'h001f,16'h0045,16'h0151,16'h0056,-16'h007c,-16'h01ce,16'h009e,16'h01b6,-16'h0024,-16'h0053,-16'h000b,16'h0103,16'h00e3,16'h0132,16'h00c4,-16'h02f5,16'h015a,16'h00bd,16'h00dd,16'h0101,-16'h0212,-16'h0432,-16'h0295,16'h0014,-16'h02e4,-16'h0175,-16'h0044,-16'h00b2,16'h00b1,16'h0036,16'h0060,-16'h0069,-16'h00e6,16'h001f,16'h00a0,-16'h0007,-16'h00e2,16'h00a7,-16'h0129,-16'h002d,16'h00ca,-16'h011e,-16'h0260,16'h014b,-16'h0052,-16'h016b,-16'h0006,16'h002b,16'h02a2,16'h000d,-16'h006d,16'h0144,16'h0048,16'h00ba,16'h010c,-16'h0029,16'h002c,-16'h012d,16'h0037,-16'h0038,16'h008b,-16'h01b3,-16'h0049,-16'h0068,16'h0095,16'h0031,16'h0088,-16'h0011,16'h0003,-16'h0144,16'h00d8,16'h016e,-16'h0029,-16'h0101,16'h002d,16'h00b7,16'h010f,16'h021a,16'h006f,-16'h0216,16'h01a9,16'h00c7,16'h0082,16'h00d8,-16'h024a,-16'h0454,-16'h0233,16'h0041,-16'h01dd,-16'h01ad,-16'h0047,-16'h005d,16'h0098,16'h0032,16'h0061,16'h0038,-16'h00b9,16'h0084,16'h00b1,16'h001c,-16'h00d4,16'h00e9,-16'h00ee,-16'h006a,16'h0060,-16'h00c2,-16'h01a8,16'h0086,16'h0025,-16'h0178,16'h0080,16'h0072,16'h0303,16'h0005,-16'h00c7,16'h00b7,16'h0065,16'h00bc,16'h00cf,-16'h0060,-16'h0040,-16'h0126,16'h000c,16'h002a,16'h0051,-16'h0386,16'h0046,-16'h0027,-16'h003c,16'h0048,16'h00d1,16'h0089,-16'h0032,16'h0003,16'h009e,16'h0159,-16'h0029,-16'h015b,16'h00d5,16'h0093,16'h016b,16'h014a,-16'h008d,-16'h022a,16'h0232,16'h00ee,16'h00a1,16'h0153,-16'h0301,-16'h034a,-16'h0114,16'h003e,-16'h01e0,-16'h0163,-16'h003f,-16'h0042,16'h00bc,16'h003e,16'h006f,16'h0041,16'h0032,16'h00a6,16'h0045,16'h00fd,-16'h00c4,16'h00b4,-16'h0136,-16'h0027,16'h008b,-16'h0075,-16'h0130,16'h0080,-16'h002e,-16'h012c,16'h00a3,16'h006f,16'h0382,16'h002a,-16'h006f,16'h0027,16'h0070,16'h0070,16'h0071,-16'h0099,-16'h0020,-16'h0100,16'h00cf,-16'h0025,16'h008b,-16'h049f,16'h00c5,-16'h0040,16'h0022,16'h0009,16'h00a7,-16'h0016,-16'h004b,16'h0074,16'h00dc,16'h01b8,-16'h0038,-16'h0168,16'h00ea,16'h0099,16'h0064,16'h017d,-16'h00a2,-16'h02ad,16'h01d7,16'h00c0,16'h00a5,16'h00fc,-16'h0386,-16'h0271,-16'h001e,-16'h0065,-16'h0216,-16'h01b3,16'h0009,16'h0046,16'h0018,16'h0068,16'h0024,16'h0094,16'h0090,16'h00cb,-16'h0083,16'h0104,-16'h00ab,16'h0052,-16'h00a9,16'h00b1,-16'h0075,-16'h001f,-16'h00cf,16'h00b8,-16'h0047,-16'h012b,16'h00bc,16'h003c,16'h02aa,16'h006b,-16'h0033,16'h0034,16'h0066,16'h009c,16'h00df,-16'h0190,16'h003a,-16'h0153,16'h010b,16'h0050,16'h006c,-16'h0499,16'h01c7,-16'h0027,16'h0002,-16'h0087,16'h0016,16'h002b,16'h0006,16'h009e,16'h00bc,16'h00be,-16'h01bf,-16'h01e9,16'h00b1,16'h002c,16'h0015,16'h0092,-16'h00ad,-16'h0290,16'h023e,16'h008c,16'h008d,16'h00d8,-16'h03a0,-16'h0105,-16'h0049,-16'h0040,-16'h017c,-16'h018a,16'h0103,-16'h0035,16'h00cb,16'h0046,16'h0016,16'h00fc,16'h0188,16'h0056,-16'h0058,16'h0163,-16'h00b7,16'h00e7,-16'h0106,16'h007b,-16'h0061,16'h001e,-16'h00e0,16'h009a,-16'h006f,-16'h01d5,16'h001a,-16'h0012,16'h0144,-16'h0015,-16'h0030,16'h0033,16'h005a,16'h0108,16'h00fc,-16'h0307,16'h0060,16'h0009,-16'h0005,16'h0000,16'h0048,-16'h038a,16'h0195,16'h004b,-16'h003b,-16'h0086,16'h0085,16'h00a4,16'h00b3,16'h00e0,16'h0019,-16'h0016,-16'h01d5,-16'h0136,16'h001c,-16'h0016,-16'h004a,16'h0036,16'h0047,-16'h0305,16'h0241,16'h0087,16'h010e,16'h00ab,-16'h0310,-16'h0068,16'h0023,-16'h0062,-16'h0154,-16'h021b,16'h016a,-16'h0025,16'h0071,16'h0100,-16'h0013,16'h013f,16'h0156,16'h00b4,-16'h0018,16'h01e8,16'h000b,16'h013e,-16'h00f5,16'h0052,-16'h0091,16'h0121,-16'h00b6,16'h0077,-16'h00c3,-16'h01ad,16'h0058,16'h0037,16'h0050,16'h001e,-16'h002d,-16'h00c3,16'h0068,16'h0174,16'h006e,-16'h040e,16'h00fb,16'h00cd,16'h0053,-16'h0056,16'h004d,-16'h0239,16'h0209,16'h008e,-16'h007c,-16'h006b,-16'h004b,16'h002c,16'h000b,16'h00a6,16'h002e,-16'h0081,-16'h01ea,-16'h00c7,16'h0064,16'h000a,-16'h00c9,16'h0059,16'h00f3,-16'h02e3,16'h02ac,16'h0088,16'h0086,16'h00be,-16'h029c,-16'h0008,16'h00d7,-16'h00d8,-16'h0174,-16'h01fd,16'h0143,-16'h00da,16'h00d5,16'h0167,16'h004f,16'h0114,16'h0132,16'h004a,16'h001c,16'h01e4,-16'h0051,16'h0188,-16'h0102,16'h0083,-16'h0076,16'h00fb,-16'h00eb,16'h0085,-16'h00d7,-16'h014b,16'h0055,-16'h0097,-16'h005c,16'h00e5,16'h0033,-16'h0136,16'h0056,16'h0133,16'h0017,-16'h02a0,16'h00bc,16'h00e2,-16'h0007,-16'h0073,16'h005c,-16'h01a9,16'h01da,16'h0058,-16'h00b7,-16'h011b,-16'h0063,16'h007e,16'h000c,16'h001a,-16'h002c,-16'h01ac,-16'h026a,-16'h00d5,-16'h006e,16'h0062,-16'h0152,16'h0085,16'h01a9,-16'h02f8,16'h0276,16'h00d6,16'h00c0,16'h0084,-16'h01d0,16'h002b,16'h0133,-16'h00f5,-16'h0199,-16'h0192,16'h01b5,-16'h010f,16'h0099,16'h016b,-16'h0075,16'h0126,16'h010d,16'h0055,16'h0019,16'h0154,16'h0081,16'h019e,-16'h012e,16'h00bc,-16'h001f,16'h007c,-16'h00d2,16'h00dc,-16'h0097,-16'h0116,-16'h0022,-16'h0030,-16'h013b,16'h005b,16'h0089,-16'h0204,16'h00b1,16'h0131,-16'h00e3,-16'h0216,16'h0159,16'h0110,16'h0021,-16'h0121,16'h00a9,-16'h0080,16'h01f4,16'h00a0,-16'h00aa,-16'h01b3,-16'h0054,16'h00b0,16'h0044,-16'h00a0,-16'h0020,-16'h0141,-16'h0142,-16'h013f,-16'h013c,16'h00b5,-16'h0197,16'h0138,16'h0187,-16'h0285,16'h0224,16'h01ab,16'h0009,16'h00e1,-16'h0177,-16'h0042,16'h0170,-16'h00f5,-16'h015a,-16'h01b6,16'h0150,-16'h0076,16'h002a,16'h00dd,-16'h0085,16'h00f0,16'h008d,16'h0014,16'h00ad,16'h011b,16'h0155,16'h00f3,-16'h0130,16'h000f,16'h00a2,16'h0092,-16'h006d,16'h0079,-16'h0011,-16'h00fe,-16'h0020,-16'h0012,-16'h0105,16'h0099,16'h00ca,-16'h02fb,16'h00af,16'h00f3,-16'h008d,-16'h0079,16'h017d,16'h005f,16'h0056,-16'h00eb,16'h002e,-16'h0076,16'h020b,16'h00e3,-16'h0031,-16'h01d1,-16'h0097,16'h011e,16'h0059,-16'h00ce,16'h0067,-16'h00bc,-16'h010a,-16'h0109,-16'h0129,16'h0176,-16'h0120,16'h01cb,16'h019e,-16'h0176,16'h01a1,16'h015d,16'h007b,16'h00bc,-16'h0082,16'h003a,16'h0132,-16'h00f6,-16'h0127,-16'h0124,16'h00f5,-16'h0085,-16'h0002,16'h0011,-16'h006a,16'h009c,16'h006b,-16'h0048,16'h00f4,16'h005f,16'h0108,16'h00a5,-16'h0138,-16'h006a,16'h0084,16'h006a,-16'h0045,16'h0051,-16'h0035,-16'h0093,16'h0097,-16'h0041,-16'h0099,16'h0033,16'h0086,-16'h02ad,16'h0068,16'h0103,-16'h0075,16'h005a,16'h012f,16'h0066,16'h003e,-16'h00bf,16'h0096,-16'h000a,16'h0150,16'h0032,-16'h009e,-16'h012b,16'h0024,16'h0029,-16'h002d,-16'h00d5,16'h009f,-16'h009c,-16'h0114,-16'h0090,-16'h00b5,16'h0123,-16'h00c2,16'h01ff,16'h00f8,-16'h00f0,16'h0173,16'h01da,16'h0073,16'h0198,-16'h00a9,-16'h0006,16'h0140,16'h0024,-16'h00fe,-16'h00e3,16'h00eb,-16'h0002,-16'h002f,16'h0033,-16'h0012,16'h00a9,16'h0088,16'h003c,16'h000c,16'h0034,16'h0132,16'h008e,-16'h00cc,16'h0015,16'h018e,16'h002f,16'h0023,16'h00db,-16'h0015,-16'h0072,16'h010a,-16'h0020,-16'h002c,16'h0054,16'h0117,-16'h02ab,-16'h004b,16'h005d,-16'h0047,16'h000c,16'h0197,16'h0045,16'h004f,-16'h00c5,16'h00c7,16'h0032,16'h017c,16'h00a0,-16'h0088,-16'h013e,16'h0054,16'h0070,-16'h001b,-16'h0095,16'h00a5,-16'h00a3,-16'h0036,-16'h00d1,-16'h0074,16'h00ab,-16'h0087,16'h01bd,16'h0023,-16'h004d,16'h00d7,16'h0233,-16'h001b,16'h01c4,-16'h0034,16'h0095,16'h0061,-16'h0038,-16'h0080,16'h0067,16'h01bb,-16'h00a5,-16'h000b,16'h0012,-16'h0014,16'h001b,16'h0051,16'h007b,-16'h004f,-16'h0045,16'h0111,16'h009d,-16'h007c,16'h0095,16'h0153,-16'h0038,16'h004a,16'h0155,16'h0045,16'h0014,16'h0118,-16'h000e,-16'h0028,-16'h0064,16'h00d8,-16'h025f,-16'h007f,16'h008c,-16'h0031,16'h004f,16'h012c,-16'h003a,16'h0053,-16'h00b2,16'h010c,-16'h0015,16'h00b5,16'h005d,-16'h0106,-16'h00e7,16'h0017,16'h005c,16'h0012,-16'h0049,16'h005e,-16'h001e,-16'h0081,-16'h0103,-16'h0086,16'h0173,-16'h006e,16'h0142,-16'h00b1,-16'h007b,16'h011c,16'h01f2,-16'h0079,16'h01e3,-16'h0011,16'h0158,16'h0031,-16'h0028,-16'h0077,16'h0114,16'h01b0,-16'h00e6,16'h0020,16'h009d,16'h0044,16'h005c,-16'h0016,-16'h0041,-16'h0085,-16'h007a,16'h00f0,16'h0087,16'h0009,16'h0052,16'h0035,-16'h007f,-16'h00a1,16'h0063,16'h0047,-16'h004a,16'h003d,16'h014e,-16'h012b,16'h003d,-16'h001e,-16'h0028,16'h0125,-16'h003b,-16'h01fa,-16'h003b,16'h018e,-16'h0043,16'h0092,-16'h0046,16'h00f0,-16'h0004,-16'h0051,16'h0083,16'h0063,-16'h0105,16'h0059,-16'h002f,16'h0070,-16'h0096,-16'h0012,-16'h00a7,-16'h0157,-16'h00c8,-16'h0091,-16'h0074,-16'h0082,16'h01b3,-16'h0088,-16'h005d,16'h00d1,-16'h0040,16'h0177,16'h0098,16'h009a,-16'h005c,-16'h00c9,16'h012e,-16'h0004,16'h007e,-16'h005f,-16'h0010,-16'h0058,-16'h00f8,16'h001c,16'h014a,-16'h01df,16'h00e1,16'h0087,16'h00de,-16'h0008,-16'h007e,-16'h00f7,-16'h00b8,-16'h0062,-16'h0080,-16'h007b,16'h00e4,16'h00c2,16'h0038,-16'h006d,16'h003d,-16'h01d8,16'h0042,16'h000a,-16'h0031,16'h011e,16'h0009,-16'h021a,16'h0074,16'h0129,16'h002d,16'h003b,16'h0067,16'h0071,-16'h000d,-16'h00b6,16'h0197,16'h0043,-16'h013a,16'h00bd,16'h0043,16'h001b,-16'h0004,16'h0047,-16'h0093,-16'h009c,-16'h0033,-16'h0013,-16'h005f,16'h0066,16'h019b,16'h009a,-16'h00fc,16'h00c8,-16'h00ee,16'h0165,16'h00a5,16'h00c7,-16'h005a,-16'h004b,16'h00ad,16'h0029,-16'h001c,-16'h00a2,-16'h00a2,-16'h00a1,16'h0009,16'h0011,16'h012e,-16'h017b,16'h002c,-16'h0033,16'h0008,-16'h004c,-16'h00ce,-16'h012e,-16'h013d,16'h0037,-16'h00aa,16'h0007,16'h011d,16'h0090,-16'h0033,-16'h000d,16'h003f,-16'h025b,16'h0068,16'h0076,-16'h007a,16'h010f,16'h0037,-16'h01b7,16'h00a9,16'h0143,-16'h0015,16'h0064,-16'h0012,16'h008f,-16'h001e,-16'h00bd,16'h029e,16'h002f,-16'h0116,16'h008c,16'h0022,16'h0063,-16'h0033,16'h001b,-16'h00bb,-16'h005c,-16'h004f,-16'h001c,-16'h00e5,-16'h0005,16'h025f,16'h0039,-16'h0124,16'h013e,-16'h00b4,16'h0138,16'h0085,16'h0113,-16'h004a,-16'h0022,16'h00b5,-16'h00bc,16'h0014,-16'h0126,-16'h019f,-16'h00b2,-16'h006a,-16'h0048,16'h00e1,-16'h008b,16'h00b6,-16'h0034,-16'h006b,-16'h0048,-16'h012b,-16'h015f,-16'h01cb,16'h008c,-16'h018a,16'h0052,16'h0121,16'h002c,-16'h00b1,-16'h00a3,16'h005c,-16'h01ee,16'h0039,16'h0038,-16'h015f,16'h0167,16'h0011,-16'h00e5,16'h0105,16'h00b4,-16'h0047,-16'h0015,16'h0019,16'h00cf,16'h0024,-16'h014c,16'h022e,16'h00ae,-16'h00b1,16'h007d,16'h000f,16'h0057,16'h000e,16'h0094,-16'h0039,-16'h005b,16'h0012,16'h00bf,-16'h017c,16'h0065,16'h02d3,16'h0015,-16'h01a6,16'h00f2,-16'h008f,16'h014f,16'h006b,16'h0130,-16'h007b,16'h007f,16'h011c,-16'h00d5,16'h0078,-16'h0124,-16'h0233,-16'h0123,-16'h003d,-16'h00ca,16'h0170,-16'h000d,16'h0060,16'h0028,-16'h012a,16'h001b,-16'h0035,-16'h0121,-16'h009d,16'h00de,-16'h01a2,16'h009a,16'h0144,-16'h0080,-16'h007f,-16'h003f,16'h0048,-16'h0178,16'h00c0,16'h0031,-16'h01a3,16'h0112,16'h0013,16'h009d,16'h00e3,-16'h006b,16'h0008,-16'h002f,-16'h0079,16'h00a9,-16'h0068,-16'h01ac,16'h01fb,16'h0059,-16'h002d,16'h0071,-16'h0080,16'h0036,-16'h0079,16'h00c3,16'h004e,16'h004e,-16'h010d,16'h00c9,-16'h0150,16'h0024,16'h025f,-16'h0043,-16'h0190,16'h00c1,16'h0016,16'h00e0,16'h00ed,16'h012a,-16'h0086,16'h0048,16'h001c,-16'h0106,16'h0158,-16'h021f,-16'h024b,-16'h00ce,-16'h005b,-16'h0090,16'h0131,16'h00ea,16'h00db,16'h004c,-16'h0152,16'h000a,-16'h00e3,-16'h010a,-16'h0025,16'h016c,-16'h02bd,16'h001c,16'h017e,-16'h008f,16'h0024,16'h0054,-16'h0043,-16'h00a2,16'h00c5,-16'h0012,-16'h022f,16'h017d,-16'h0041,16'h007a,16'h0056,-16'h019b,-16'h006e,16'h0074,16'h0015,16'h0122,16'h0075,-16'h0107,16'h00a9,16'h0016,-16'h0018,16'h00d5,-16'h0041,16'h0061,-16'h0027,16'h00d2,16'h00cc,16'h006a,-16'h0127,16'h0081,-16'h0199,16'h0025,16'h027a,-16'h0082,-16'h019b,16'h0128,16'h008d,16'h00fe,16'h00ac,16'h0132,-16'h00b1,16'h0089,-16'h001e,-16'h013f,16'h011a,-16'h023c,-16'h0104,-16'h0129,16'h0031,-16'h0056,16'h0102,16'h00e5,16'h00de,16'h00cb,-16'h00fb,16'h0047,-16'h00bc,-16'h0134,16'h0026,16'h017b,-16'h02c7,16'h004e,16'h01d4,-16'h001b,-16'h006d,-16'h0023,-16'h00cf,-16'h0097,16'h0045,-16'h00b8,-16'h026a,16'h0140,16'h0048,16'h010c,-16'h000a,-16'h01bf,-16'h003f,16'h004b,-16'h0016,16'h0051,16'h00a3,-16'h0145,-16'h0153,16'h0079,16'h000a,16'h0159,16'h000d,-16'h001a,16'h0048,-16'h000a,16'h013c,16'h00d1,-16'h0185,16'h00cb,-16'h0042,16'h0094,16'h0218,-16'h007b,-16'h01b5,16'h00c8,16'h00e8,-16'h0018,16'h0031,16'h00d7,-16'h00f7,16'h0013,-16'h0088,-16'h0253,16'h00a4,-16'h02a2,-16'h0015,-16'h0130,16'h003a,16'h000d,16'h0131,16'h00ae,-16'h000b,16'h00e4,16'h001a,16'h002b,-16'h008d,-16'h008c,16'h0012,16'h0167,-16'h0261,16'h0118,16'h01ef,16'h0004,-16'h001b,-16'h009e,-16'h0109,-16'h00af,-16'h0059,-16'h00cc,-16'h020f,16'h012b,-16'h001b,16'h00d0,16'h003c,-16'h01a4,-16'h00b2,16'h002e,16'h004b,16'h0062,16'h008a,-16'h010f,-16'h02f0,16'h0030,-16'h0016,16'h00e1,16'h0044,16'h0020,16'h0064,16'h005a,16'h0088,16'h00a6,-16'h0195,16'h0017,16'h0025,16'h003d,16'h01c6,-16'h004b,-16'h0221,16'h014e,16'h0036,16'h0017,16'h0032,16'h0112,-16'h013f,16'h0001,-16'h0005,-16'h02d7,16'h0013,-16'h0218,16'h0014,-16'h00ea,16'h012d,-16'h0020,16'h0130,16'h0144,16'h0014,16'h00ed,16'h0013,16'h0021,-16'h0044,-16'h0073,16'h0045,16'h012c,-16'h01ca,16'h00f7,16'h024e,16'h0037,-16'h0019,-16'h0022,-16'h00c6,16'h004c,-16'h007c,-16'h010c,-16'h01ce,16'h0088,-16'h0052,16'h00ba,16'h001c,-16'h0090,-16'h0048,16'h0032,16'h000e,16'h001c,16'h00ab,-16'h0158,-16'h0391,16'h0100,-16'h0067,16'h00bb,16'h005c,-16'h009b,16'h0028,-16'h0015,16'h01ae,-16'h0017,-16'h01a7,16'h0012,16'h0074,-16'h00c6,16'h01bb,-16'h00eb,-16'h01ff,16'h012e,16'h008e,-16'h000f,16'h009a,16'h0064,-16'h01d3,-16'h00c9,-16'h0078,-16'h0288,-16'h0082,-16'h01a5,16'h0013,-16'h0070,16'h00e7,16'h0080,16'h00c5,16'h00f0,16'h001e,16'h010a,16'h0083,16'h005c,16'h0014,-16'h0065,16'h0060,16'h0133,-16'h0152,16'h0080,16'h0282,16'h0000,-16'h000e,-16'h005a,-16'h0023,16'h002e,-16'h004d,-16'h00fa,-16'h00fa,-16'h0029,-16'h003c,-16'h004d,-16'h0003,-16'h00ea,-16'h000a,-16'h003e,-16'h0026,16'h004d,16'h00bd,-16'h00d0,-16'h0492,16'h0080,-16'h0030,16'h0089,16'h009e,-16'h009a,16'h00b2,-16'h007b,16'h0146,16'h0038,-16'h0171,16'h0000,16'h011f,-16'h00c7,16'h01e3,-16'h004d,-16'h026b,16'h0105,16'h0005,-16'h006f,16'h0101,-16'h0027,-16'h01d0,-16'h0145,-16'h00bb,-16'h01e1,-16'h0065,-16'h0097,-16'h0041,-16'h0062,16'h0070,16'h002d,16'h006a,16'h00da,-16'h008b,16'h0052,16'h001d,16'h0035,16'h0084,-16'h009f,16'h0059,16'h0108,-16'h00d2,16'h001c,16'h0247,-16'h000f,-16'h000b,-16'h0068,-16'h0086,16'h00ef,16'h002b,-16'h00cd,-16'h008c,-16'h009b,-16'h0046,-16'h0074,16'h004c,-16'h0113,16'h0028,16'h002f,16'h000c,16'h0000,16'h00a3,-16'h0136,-16'h0404,16'h004d,-16'h0004,16'h005f,16'h00ea,-16'h0006,16'h004d,-16'h00e9,16'h01a2,-16'h0013,-16'h00f6,-16'h0049,16'h0150,-16'h00df,16'h0227,16'h002c,-16'h0269,16'h0174,-16'h0036,16'h000e,16'h00a8,-16'h0078,-16'h0261,-16'h01c0,-16'h005e,-16'h01fd,-16'h00b2,-16'h0019,-16'h0025,-16'h0056,16'h0096,-16'h0005,-16'h0022,16'h001b,-16'h004f,16'h00d2,-16'h00a0,-16'h000a,16'h0024,-16'h0044,-16'h00cc,16'h001b,-16'h011d,-16'h0064,16'h0206,-16'h006b,16'h005c,-16'h0056,16'h0004,16'h00ec,16'h003a,-16'h00d8,-16'h0056,-16'h00bb,-16'h0011,-16'h0101,16'h006a,-16'h0139,16'h000c,-16'h0071,-16'h007d,-16'h0039,16'h0106,-16'h00da,-16'h033d,16'h0077,16'h0027,16'h006a,16'h014a,-16'h0025,16'h003d,-16'h00a0,16'h0121,-16'h001c,-16'h011a,-16'h005d,16'h0178,-16'h0011,16'h0226,16'h001d,-16'h0270,16'h0146,-16'h001b,16'h0047,16'h0074,-16'h0088,-16'h0321,-16'h027f,-16'h005f,-16'h0213,-16'h00dd,16'h001c,-16'h0021,16'h0024,16'h0074,16'h003f,-16'h001d,-16'h00c1,-16'h00d7,16'h00bd,-16'h00b8,-16'h0023,16'h00c1,-16'h00a6,-16'h001e,16'h006c,-16'h00d6,-16'h00fa,16'h0154,-16'h0005,16'h0068,-16'h0021,16'h0059,16'h01d1,16'h0081,-16'h0055,-16'h0078,-16'h0086,16'h0044,16'h0002,16'h0093,-16'h00bb,-16'h0011,-16'h005b,-16'h0087,16'h0023,16'h012e,-16'h011f,-16'h0253,16'h002e,-16'h0014,16'h0023,16'h00a6,-16'h005d,-16'h0038,-16'h00ef,16'h00f1,16'h0015,-16'h00a8,-16'h0022,16'h016a,-16'h0017,16'h01c1,16'h003b,-16'h027a,16'h00fe,-16'h002f,16'h0023,16'h0080,-16'h006d,-16'h046e,-16'h039d,-16'h009b,-16'h0253,-16'h00ce,-16'h004a,-16'h0022,16'h0051,16'h008a,16'h002f,-16'h0071,-16'h01ff,-16'h0062,16'h008b,-16'h0070,16'h0023,-16'h002a,-16'h0087,-16'h003a,16'h00d4,16'h0012,-16'h0175,16'h018c,16'h003e,16'h0036,-16'h0024,16'h0071,16'h021b,16'h005e,-16'h0027,16'h0075,-16'h00af,16'h0069,16'h009a,16'h00e1,-16'h0067,-16'h001b,-16'h00bd,-16'h004c,16'h003b,16'h0114,-16'h016b,-16'h0123,16'h0005,16'h008e,16'h0066,16'h00e6,-16'h009c,-16'h003e,-16'h0026,16'h00bd,16'h0038,-16'h007e,-16'h001b,16'h0153,-16'h0002,16'h01ef,16'h00a6,-16'h028f,16'h016c,16'h005b,-16'h0030,16'h0027,-16'h0071,-16'h040b,-16'h0365,-16'h0024,-16'h0281,-16'h0142,-16'h000c,-16'h0089,16'h005e,16'h00b7,16'h00f6,-16'h006c,-16'h01cb,-16'h0023,16'h013e,-16'h0077,-16'h0010,-16'h0024,-16'h00de,-16'h0004,16'h0030,16'h0024,-16'h0252,16'h015b,16'h0055,16'h0063,16'h0039,16'h00ba,16'h01bb,16'h0044,-16'h000c,16'h00e1,-16'h009a,16'h000b,16'h0187,16'h0051,-16'h000d,-16'h0007,-16'h00a5,16'h001b,16'h008b,16'h010a,-16'h0071,-16'h0062,-16'h002a,16'h0032,16'h00a7,16'h003d,-16'h007b,-16'h00d9,16'h0008,16'h00ab,16'h000c,-16'h0093,-16'h0037,16'h0092,16'h002c,16'h0223,16'h00ed,-16'h022e,16'h0151,16'h00b1,-16'h004d,16'h00c2,-16'h0049,-16'h03a8,-16'h036b,-16'h0009,-16'h027f,-16'h01fe,-16'h0065,-16'h003c,16'h00a4,16'h008f,16'h00cb,-16'h009c,-16'h012e,16'h0014,16'h00ad,-16'h0032,16'h0000,16'h0023,-16'h00de,-16'h0072,-16'h0009,16'h0090,-16'h01aa,16'h0190,-16'h0062,-16'h0048,-16'h0039,16'h0075,16'h01f5,16'h0028,16'h0028,16'h011f,-16'h00c9,16'h0099,16'h014f,16'h0046,16'h0028,-16'h005d,-16'h00d1,-16'h0025,16'h004d,16'h002d,-16'h000f,16'h0014,-16'h0029,16'h004f,16'h0057,-16'h002e,-16'h0045,-16'h0122,16'h003c,16'h0107,16'h0017,-16'h005c,16'h001b,16'h000b,16'h00c5,16'h01d2,16'h0119,-16'h0216,16'h0204,16'h0056,16'h003d,16'h00f5,-16'h00c9,-16'h0313,-16'h034e,16'h0081,-16'h025a,-16'h01a7,-16'h0046,16'h000e,16'h0059,16'h0016,16'h011b,16'h003c,-16'h005e,16'h004b,16'h0079,16'h0063,-16'h0050,-16'h000d,-16'h00ee,-16'h0063,-16'h003d,16'h001d,-16'h0072,16'h0174,-16'h0039,-16'h00dc,16'h000d,16'h0016,16'h0242,-16'h0011,16'h008b,16'h0137,-16'h00ae,16'h002a,16'h0090,16'h00a5,-16'h0011,-16'h0098,-16'h0024,-16'h003b,-16'h0004,-16'h0060,16'h0041,16'h00cc,-16'h0069,16'h0021,16'h00bb,-16'h002d,16'h0036,-16'h00e4,16'h0011,16'h0133,-16'h0031,-16'h004e,16'h0083,16'h0061,16'h0139,16'h021f,16'h0109,-16'h0192,16'h01dc,16'h00af,-16'h0096,16'h0072,-16'h012e,-16'h0347,-16'h033e,16'h0056,-16'h01e6,-16'h015d,16'h000d,16'h0065,16'h007b,-16'h0025,16'h0165,16'h0072,-16'h006e,16'h0086,-16'h0021,16'h0071,-16'h00e2,16'h00c4,-16'h002f,-16'h0030,16'h001b,-16'h0021,-16'h0034,16'h0114,16'h003f,-16'h01e2,16'h002e,-16'h000a,16'h027a,-16'h0045,16'h003f,16'h0118,16'h001b,-16'h00a7,-16'h001d,16'h011a,-16'h0005,-16'h008d,-16'h004a,-16'h0039,16'h0027,-16'h02b1,16'h00e2,16'h00c0,-16'h0134,-16'h0033,16'h007a,-16'h00ac,-16'h006b,-16'h0063,16'h0034,16'h0104,-16'h0013,-16'h0116,16'h00c3,16'h0082,16'h010a,16'h01df,16'h0018,-16'h01e9,16'h01d3,16'h00bd,-16'h006a,16'h0016,-16'h022f,-16'h0280,-16'h0265,16'h004c,-16'h017e,-16'h01c1,16'h0013,16'h0004,16'h002e,-16'h003e,16'h010b,16'h00be,16'h007b,16'h005a,16'h0006,16'h006b,-16'h00e0,16'h0007,-16'h00a9,-16'h0062,16'h0016,16'h000c,16'h0011,16'h00c7,16'h0027,-16'h0116,16'h0000,16'h0053,16'h0234,-16'h0081,-16'h0021,16'h0083,16'h001c,-16'h0056,16'h001a,-16'h005e,16'h0063,-16'h00f5,16'h004c,16'h0097,-16'h001e,-16'h049d,16'h0128,16'h006c,-16'h00df,-16'h006a,16'h0087,-16'h008a,-16'h002c,-16'h0008,16'h00a7,16'h00e2,-16'h00c4,-16'h01a1,16'h0095,16'h0041,16'h0121,16'h0160,-16'h00bd,-16'h0178,16'h01fa,16'h0082,16'h000a,16'h0059,-16'h02ce,-16'h0166,-16'h0140,16'h00d1,-16'h01c6,-16'h01b4,16'h000f,16'h004a,16'h00db,-16'h0003,16'h0123,16'h0090,16'h013a,16'h00db,-16'h00f8,16'h00d5,-16'h00d0,-16'h000d,-16'h00b0,16'h008d,-16'h0004,16'h000a,-16'h0015,16'h0099,-16'h0008,-16'h0133,-16'h001d,-16'h0009,16'h016c,-16'h006b,-16'h0010,16'h005d,16'h0071,16'h0036,16'h0050,-16'h0101,16'h006f,-16'h011f,16'h005d,16'h001c,16'h006f,-16'h0555,16'h0124,-16'h000a,-16'h007b,-16'h00a1,16'h0002,-16'h0084,-16'h0031,16'h00be,16'h00bc,16'h002c,-16'h00f0,-16'h01c6,16'h0070,-16'h006c,16'h0097,16'h00df,-16'h009c,-16'h0140,16'h0234,16'h008a,16'h00b1,16'h0074,-16'h036e,-16'h007a,-16'h0118,16'h0056,-16'h01d1,-16'h01ab,16'h0000,16'h005f,16'h00c1,-16'h000d,16'h00ea,16'h00e7,16'h0133,16'h0039,-16'h00c1,16'h00e3,-16'h007b,16'h002b,-16'h00a8,16'h00c0,-16'h0004,16'h005c,-16'h0062,16'h008c,-16'h000a,-16'h0126,-16'h0003,16'h0048,16'h008c,16'h0006,-16'h0023,-16'h0018,16'h009e,16'h0050,16'h0078,-16'h02ec,16'h00a7,-16'h00b9,-16'h002f,16'h004e,16'h0009,-16'h03c8,16'h0136,16'h0052,-16'h005a,-16'h0016,16'h0008,16'h0044,16'h006a,16'h0170,16'h004f,-16'h00ee,-16'h0188,-16'h010d,-16'h0037,-16'h00bb,16'h001e,16'h00a4,16'h0001,-16'h01b6,16'h02aa,16'h001d,16'h00cc,16'h0009,-16'h038a,16'h004d,-16'h0090,16'h000f,-16'h01f7,-16'h01a5,16'h00ea,16'h0029,16'h010b,16'h008a,16'h0022,16'h0074,16'h0112,16'h0097,-16'h00c7,16'h012c,-16'h0040,16'h003e,-16'h005c,16'h0132,16'h0006,16'h00a7,-16'h011a,16'h005b,16'h0028,-16'h00bd,-16'h001b,-16'h0026,-16'h007e,16'h0086,-16'h0070,-16'h0040,16'h00e0,16'h00a0,16'h0010,-16'h0534,16'h00e8,-16'h0019,16'h0042,16'h001f,16'h0103,-16'h01e4,16'h0172,16'h003e,16'h005b,-16'h0083,-16'h004e,16'h0066,16'h004c,16'h00cc,-16'h0082,-16'h01dd,-16'h014f,-16'h009d,-16'h0060,-16'h0054,-16'h00ed,16'h0040,16'h008a,-16'h01b4,16'h021a,16'h00ee,16'h00d9,-16'h006e,-16'h0361,16'h009c,-16'h0027,16'h0059,-16'h0111,-16'h01ff,16'h006f,16'h000d,16'h008f,16'h0114,-16'h000a,16'h00f8,16'h00bd,16'h00f7,-16'h003d,16'h01e0,16'h0072,16'h0009,-16'h0048,16'h0137,-16'h0041,16'h0146,-16'h0064,16'h007d,16'h00a9,-16'h0068,16'h0006,-16'h001c,-16'h011e,16'h0070,-16'h0067,-16'h0130,16'h0148,16'h00bc,-16'h00a5,-16'h03d5,16'h00ac,16'h00c0,16'h006e,-16'h0057,16'h0155,-16'h018c,16'h010c,16'h006a,-16'h00ab,-16'h00af,-16'h0005,16'h00c5,16'h0037,16'h0059,-16'h00e8,-16'h0221,-16'h014d,-16'h0096,-16'h0068,-16'h0003,-16'h008e,16'h007c,16'h022b,-16'h0159,16'h0212,16'h009a,16'h00dd,-16'h005a,-16'h027c,16'h00b4,16'h0040,-16'h0094,-16'h016c,-16'h00f2,16'h00dd,-16'h008a,16'h00bf,16'h0114,-16'h0043,16'h00fb,16'h00f7,16'h0166,16'h0029,16'h0161,16'h00ef,16'h0028,-16'h00c2,16'h008c,-16'h0079,16'h0138,16'h002e,16'h00bd,16'h0075,-16'h0098,-16'h001c,-16'h002d,-16'h018f,16'h0027,-16'h0083,-16'h023b,16'h0133,16'h00f3,-16'h00bc,-16'h0281,16'h0120,16'h00fd,16'h002d,-16'h00b6,16'h0060,-16'h00b4,16'h00e2,16'h00a9,-16'h00cd,-16'h0131,-16'h0027,16'h00d8,16'h0017,16'h0021,-16'h0103,-16'h01ec,-16'h010a,-16'h0106,16'h0009,16'h000e,-16'h00a7,16'h0118,16'h023f,-16'h0129,16'h0262,16'h0107,16'h00de,-16'h00a4,-16'h018e,16'h010e,16'h00c8,-16'h00e1,-16'h0193,-16'h00da,16'h00de,-16'h0054,16'h00a2,16'h006f,-16'h007e,16'h0139,16'h0089,16'h00db,16'h00e6,16'h017a,16'h0155,16'h0052,-16'h0113,16'h00be,16'h0060,16'h00eb,16'h007c,16'h00ad,16'h005d,-16'h0076,-16'h00b1,-16'h007c,-16'h0172,-16'h0007,16'h006a,-16'h033a,16'h0148,16'h00e3,-16'h00d3,-16'h0100,16'h00a9,16'h00d6,-16'h0075,-16'h00d4,16'h002d,-16'h0027,16'h010d,16'h0062,-16'h0136,-16'h0148,-16'h0063,16'h006f,-16'h0033,16'h0040,-16'h006d,-16'h016c,-16'h0122,-16'h0157,-16'h009d,16'h0036,-16'h013d,16'h01cc,16'h0237,-16'h00dc,16'h021c,16'h00cb,16'h0090,16'h0012,-16'h00e4,16'h010d,16'h0100,-16'h0104,-16'h01e3,-16'h00a2,16'h0134,-16'h00b4,16'h0015,-16'h0001,-16'h0109,16'h0047,16'h006f,16'h004d,16'h01ac,16'h008f,16'h01ca,16'h0022,-16'h00ea,16'h0085,16'h0089,16'h00ea,16'h0029,16'h0079,-16'h0003,-16'h0036,-16'h0041,-16'h0030,-16'h00b9,16'h00b9,16'h0096,-16'h02cc,16'h0092,16'h00f9,-16'h00ac,16'h006c,16'h0118,16'h008b,-16'h009f,-16'h00ec,16'h0067,16'h0037,16'h00a4,16'h0029,-16'h00be,-16'h016e,-16'h002c,16'h005b,16'h0079,-16'h00ef,16'h00c0,-16'h0115,-16'h00a8,-16'h0122,-16'h0056,16'h008d,-16'h00a1,16'h01d9,16'h01e2,-16'h0030,16'h0186,16'h012e,16'h008c,16'h00b1,-16'h0039,16'h00ec,16'h0105,-16'h0012,-16'h0160,-16'h00c1,16'h016f,-16'h0009,16'h0036,-16'h001b,-16'h0026,-16'h002e,16'h00c9,16'h0014,16'h0124,16'h005c,16'h0135,16'h009d,-16'h006c,-16'h0009,16'h00bc,16'h0024,16'h008d,16'h0054,16'h001b,16'h0017,16'h00c0,16'h000a,-16'h003c,16'h00a1,16'h00cc,-16'h02f6,16'h00c4,16'h00b6,-16'h001f,16'h00f0,16'h016f,16'h003e,-16'h0001,-16'h004e,16'h0090,16'h000b,16'h009c,16'h0015,-16'h00a8,-16'h012e,16'h001d,16'h001c,-16'h004c,-16'h00b1,16'h012b,-16'h007d,-16'h00a0,-16'h0169,-16'h00c5,16'h006e,-16'h00df,16'h021d,16'h011f,-16'h0008,16'h011d,16'h0219,16'h003d,16'h015a,-16'h0001,16'h00e4,16'h00c7,-16'h0025,-16'h0131,-16'h0052,16'h018f,-16'h0069,16'h005d,16'h0006,-16'h0088,16'h004b,16'h0002,16'h002c,16'h000e,-16'h005c,16'h015e,16'h00f6,-16'h0038,16'h003d,16'h00d9,16'h0098,16'h0080,16'h00a2,16'h00ac,-16'h006c,16'h0129,-16'h0063,-16'h00c2,16'h0028,16'h00ce,-16'h0250,-16'h0078,16'h0073,-16'h003e,16'h00b4,16'h01a9,16'h0066,16'h0057,-16'h0039,16'h008f,-16'h0015,16'h0093,16'h0049,-16'h00b9,-16'h00f0,16'h0052,16'h004f,-16'h0035,-16'h00a5,16'h00bc,-16'h004b,-16'h00ce,-16'h011a,-16'h0008,16'h003b,-16'h0039,16'h01b0,-16'h0033,16'h0009,16'h00c5,16'h01f5,16'h0034,16'h0171,-16'h0036,16'h00f6,16'h00e9,-16'h0063,-16'h006e,16'h0059,16'h0186,-16'h00e1,16'h0044,16'h008a,-16'h005b,16'h00b8,-16'h0009,16'h0075,-16'h005d,-16'h0086,16'h017e,16'h00cf,16'h0017,16'h0047,16'h0020,-16'h003d,-16'h0140,16'h00a3,16'h0032,-16'h004f,16'h0074,16'h00f5,-16'h0185,16'h0007,16'h000a,16'h0098,16'h0074,-16'h0051,-16'h0201,16'h00a3,16'h0183,16'h001f,16'h0039,16'h004c,16'h0089,-16'h0087,-16'h0014,16'h0139,16'h00c3,-16'h015f,16'h00e4,-16'h0035,16'h003f,16'h0030,16'h0019,-16'h00fe,-16'h0127,-16'h008f,-16'h00c9,-16'h003d,16'h0021,16'h0163,16'h00b9,-16'h003a,16'h010a,-16'h00ca,16'h0190,16'h00bc,16'h00a1,-16'h00a1,-16'h00cf,16'h00f2,16'h0020,16'h0099,-16'h00cf,-16'h0002,-16'h00e9,-16'h00c7,16'h0054,16'h0136,-16'h018f,16'h00c3,-16'h0062,16'h00ed,-16'h002f,-16'h0057,-16'h00da,-16'h00c2,-16'h00bc,-16'h00a5,-16'h005a,16'h00f3,16'h00a9,-16'h0031,-16'h0033,16'h00af,-16'h025a,16'h011e,-16'h0010,-16'h0025,16'h00e3,-16'h000c,-16'h015b,16'h013b,16'h0166,16'h006f,16'h007b,-16'h0035,16'h0045,-16'h0079,-16'h007e,16'h02c0,16'h00f9,-16'h0115,16'h00c1,16'h0002,16'h0015,16'h0085,16'h005b,-16'h011c,-16'h0050,-16'h0095,16'h0028,16'h000b,16'h00a7,16'h01b6,16'h00cd,-16'h00ac,16'h00ca,-16'h00b0,16'h0174,16'h008b,16'h00cc,-16'h00bb,-16'h00bf,16'h008b,-16'h0013,-16'h0016,-16'h013a,-16'h0170,-16'h00df,-16'h0005,-16'h00b9,16'h016b,-16'h00a5,16'h0074,-16'h0006,-16'h0046,-16'h009f,-16'h00d9,-16'h0103,-16'h00d0,-16'h000d,-16'h00ab,-16'h0033,16'h01a9,-16'h0047,-16'h00b6,-16'h009b,16'h00e9,-16'h0278,16'h00d4,16'h00b2,-16'h00b1,16'h00e4,16'h0027,-16'h0103,16'h0108,16'h0169,16'h009f,16'h0036,-16'h0042,16'h007c,-16'h00c5,-16'h012a,16'h02c4,16'h0077,-16'h00ef,16'h00f6,-16'h000d,-16'h0026,16'h0071,16'h006b,-16'h00f7,-16'h0030,-16'h002f,16'h005a,-16'h00db,16'h0050,16'h022b,16'h0011,-16'h00ff,16'h0147,-16'h0094,16'h01e6,16'h00c9,16'h009c,-16'h00cb,-16'h001e,16'h0165,-16'h0132,16'h00a3,-16'h01a5,-16'h01a6,-16'h0139,-16'h0068,-16'h00b5,16'h0150,-16'h0083,16'h00a7,16'h0047,-16'h005f,-16'h0082,-16'h0061,-16'h00fb,-16'h00af,16'h00da,-16'h0173,-16'h0010,16'h01b2,-16'h00c1,-16'h00cc,16'h0013,16'h00fb,-16'h01ff,16'h006e,16'h0090,-16'h015b,16'h019d,16'h0062,16'h004a,16'h00d0,16'h0081,16'h0024,16'h0042,-16'h008a,16'h00b9,-16'h008c,-16'h0112,16'h027d,16'h0069,-16'h005c,16'h00ed,16'h000d,-16'h004f,-16'h004f,16'h003a,-16'h0026,-16'h000a,-16'h00cc,16'h00b4,-16'h014c,16'h005a,16'h0218,16'h003b,-16'h009c,16'h010e,-16'h00a2,16'h0135,16'h00f1,16'h007c,-16'h00ce,16'h0057,16'h00a5,-16'h00b7,16'h011a,-16'h0239,-16'h027d,-16'h00e8,-16'h0068,-16'h00fd,16'h012e,16'h0020,16'h00d5,16'h002b,-16'h008d,16'h0006,-16'h000c,-16'h0085,-16'h0034,16'h0101,-16'h0296,16'h000f,16'h028b,-16'h0101,-16'h0088,16'h004e,16'h0061,-16'h01a1,16'h00a1,16'h003d,-16'h0267,16'h015d,16'h0047,16'h003e,16'h00d9,-16'h008d,16'h005a,16'h0029,-16'h0057,16'h00c6,-16'h0037,-16'h012f,16'h0181,16'h0066,-16'h0001,16'h00a9,-16'h0099,-16'h0007,-16'h0002,16'h003f,-16'h0038,16'h002e,-16'h0145,16'h005f,-16'h0115,16'h0050,16'h0209,-16'h0044,-16'h0053,16'h011d,-16'h001f,16'h00bd,16'h008e,16'h010b,-16'h00db,16'h0081,16'h004f,-16'h0105,16'h012d,-16'h02f1,-16'h01ff,-16'h014f,-16'h0023,-16'h008b,16'h0118,16'h007e,16'h00c7,16'h005c,16'h0032,-16'h009d,-16'h00a0,-16'h0058,-16'h0069,16'h00eb,-16'h02e5,16'h0030,16'h028c,-16'h00ea,-16'h0010,16'h0041,16'h005a,-16'h00a6,16'h003d,-16'h002e,-16'h02d2,16'h0160,16'h0004,16'h0101,16'h0051,-16'h01d1,16'h0065,-16'h000a,-16'h0011,16'h00dd,16'h001f,-16'h0133,-16'h003b,16'h0044,-16'h0047,16'h00b4,-16'h0088,-16'h001d,16'h0000,16'h0061,16'h00b9,16'h0046,-16'h01c9,16'h00a6,-16'h00f4,16'h00b5,16'h0245,-16'h007a,-16'h0005,16'h00ab,16'h009e,16'h00cd,16'h00c2,16'h0135,-16'h00a6,16'h0015,-16'h001b,-16'h0175,16'h0171,-16'h031b,-16'h0079,-16'h018a,16'h007c,-16'h0074,16'h01b6,16'h00ed,16'h00ad,16'h0074,-16'h002d,16'h0035,-16'h001d,-16'h0073,-16'h002f,16'h0172,-16'h0310,16'h0102,16'h024b,-16'h0055,-16'h003e,16'h00bc,-16'h0045,-16'h0072,-16'h002d,-16'h00af,-16'h02bb,16'h012c,16'h002d,16'h0092,16'h0078,-16'h019e,16'h001c,-16'h004e,-16'h0088,16'h009c,16'h0033,-16'h0161,-16'h0207,16'h009c,-16'h007e,16'h00ec,-16'h0083,-16'h0053,-16'h0017,16'h0001,16'h0104,16'h0092,-16'h0194,-16'h000e,16'h0001,-16'h000c,16'h0227,-16'h00f6,-16'h002e,16'h0148,16'h00a7,-16'h0037,16'h004d,16'h012c,-16'h00e6,-16'h002c,-16'h006b,-16'h0217,16'h00be,-16'h02d0,-16'h0017,-16'h0172,16'h00c3,16'h0015,16'h0149,16'h0117,16'h0089,16'h00fe,-16'h002d,16'h0013,-16'h000b,-16'h0099,16'h0004,16'h0156,-16'h01b0,16'h0124,16'h028a,-16'h0028,-16'h003b,16'h001f,-16'h00b3,16'h0002,-16'h002a,-16'h0083,-16'h0254,16'h00bd,-16'h007c,16'h001b,-16'h000e,-16'h0102,16'h0044,-16'h0034,-16'h006b,16'h00a5,16'h0036,-16'h01da,-16'h0435,16'h0084,-16'h0013,16'h00b0,-16'h0020,-16'h002a,16'h0047,16'h0098,16'h00eb,16'h0025,-16'h0132,16'h0016,16'h0085,16'h003f,16'h027c,-16'h00e8,-16'h0051,16'h013d,16'h008c,16'h0080,16'h00cf,16'h00a2,-16'h0166,-16'h0062,16'h0009,-16'h0273,-16'h001c,-16'h0122,-16'h008e,-16'h019a,16'h0128,16'h002b,16'h00cd,16'h0103,16'h004c,16'h00e4,16'h0011,-16'h0001,16'h004a,-16'h007b,16'h0015,16'h017d,-16'h0105,16'h010d,16'h0280,-16'h0056,-16'h004c,-16'h0014,-16'h008e,16'h003b,-16'h0055,-16'h011f,-16'h01aa,16'h00b7,-16'h0046,-16'h002f,-16'h0019,-16'h0195,-16'h000b,16'h000a,-16'h0016,16'h0099,16'h0030,-16'h017d,-16'h04b3,16'h010f,16'h002e,16'h0071,-16'h0051,-16'h003f,16'h0015,-16'h0013,16'h017f,-16'h000e,-16'h00ef,-16'h003c,16'h0101,-16'h00b9,16'h02cb,-16'h00c9,-16'h003c,16'h0156,16'h003c,16'h0041,16'h00ee,16'h0039,-16'h0195,-16'h003c,-16'h00e8,-16'h027f,-16'h006a,-16'h00a8,-16'h004b,-16'h0155,16'h0097,16'h004d,16'h006b,16'h0185,16'h0003,16'h00c9,16'h0004,16'h00be,16'h0015,-16'h00df,-16'h006f,16'h0065,-16'h0056,16'h0019,16'h0285,-16'h0081,-16'h0015,-16'h009e,-16'h00f4,16'h001b,-16'h0036,-16'h00c8,-16'h0165,16'h0009,16'h003b,-16'h0038,16'h009d,-16'h0191,-16'h0029,-16'h002c,16'h002a,-16'h0020,16'h00ba,-16'h01a1,-16'h0473,16'h0043,-16'h0023,16'h002b,-16'h0003,-16'h0058,16'h003c,-16'h0063,16'h01a5,-16'h0006,-16'h008c,16'h0045,16'h014b,-16'h0059,16'h0271,-16'h0072,-16'h006a,16'h0179,16'h0027,16'h0062,16'h0048,-16'h000f,-16'h026d,-16'h00b9,-16'h00c3,-16'h024c,-16'h009e,16'h004f,-16'h0057,-16'h0143,16'h006f,16'h000a,16'h0036,16'h00d0,16'h0009,16'h007b,-16'h0054,16'h0012,-16'h0017,-16'h00e0,-16'h008d,16'h0058,-16'h0021,-16'h0002,16'h0299,-16'h0055,-16'h0002,-16'h0055,-16'h0030,16'h00ad,16'h0001,-16'h00d5,-16'h00d6,-16'h006c,-16'h001f,-16'h005d,16'h0052,-16'h0154,-16'h0079,-16'h0053,-16'h0064,16'h0048,16'h00d2,-16'h0115,-16'h037f,16'h0082,16'h0014,16'h006f,16'h002e,-16'h0005,16'h0065,-16'h00a7,16'h0122,-16'h0064,-16'h008b,-16'h0027,16'h01b2,-16'h000c,16'h024f,16'h0025,-16'h0076,16'h0177,16'h001c,16'h002d,16'h00d7,-16'h0055,-16'h038c,-16'h00ef,-16'h007f,-16'h028f,-16'h00a4,16'h0065,-16'h0071,-16'h00b2,16'h0065,-16'h003d,16'h001a,-16'h00ab,16'h0017,16'h00ad,-16'h008d,16'h0078,-16'h0019,-16'h0133,-16'h000b,16'h000c,16'h00ad,-16'h00d0,16'h01fe,-16'h004a,16'h00f6,-16'h005e,16'h0033,16'h0154,16'h0042,-16'h00c9,-16'h00f7,-16'h0063,-16'h000e,-16'h0098,16'h0019,-16'h0105,-16'h0086,-16'h00ab,16'h0012,16'h0020,16'h0147,-16'h0128,-16'h0263,16'h0082,-16'h0079,16'h004e,16'h00db,-16'h0042,16'h0021,-16'h00e6,16'h012c,-16'h0069,-16'h007d,16'h000c,16'h0141,16'h0077,16'h026c,-16'h0013,-16'h0067,16'h019d,16'h0051,16'h0032,16'h0086,-16'h0036,-16'h0474,-16'h01ad,-16'h00a8,-16'h0262,-16'h00c0,-16'h0089,-16'h003f,-16'h00a7,16'h005f,16'h0072,16'h001e,-16'h0153,-16'h0061,16'h00a0,-16'h004f,16'h000d,-16'h0034,-16'h00b2,-16'h001e,16'h0075,16'h0049,-16'h00de,16'h01d1,16'h0025,16'h00d9,-16'h008f,16'h0031,16'h0191,16'h0076,16'h003a,-16'h00e6,-16'h012b,-16'h0014,16'h0094,-16'h0011,-16'h0075,16'h000e,-16'h002f,-16'h002c,16'h0042,16'h013a,-16'h01ac,-16'h00e6,16'h002e,16'h001d,-16'h0042,16'h00e0,-16'h0027,-16'h003f,-16'h0058,16'h00a9,-16'h0050,-16'h0017,16'h0053,16'h00aa,-16'h0019,16'h0271,16'h00a4,-16'h003d,16'h0137,16'h0026,-16'h0013,16'h00db,16'h000a,-16'h04b3,-16'h0287,-16'h0047,-16'h0281,-16'h0105,16'h005c,-16'h0072,-16'h006f,16'h0036,16'h003c,-16'h0067,-16'h01c6,-16'h0060,16'h0116,-16'h002d,-16'h0029,16'h0016,-16'h0081,-16'h0002,16'h0033,16'h0048,-16'h0138,16'h0225,-16'h0006,16'h00ec,-16'h0080,16'h0026,16'h0227,16'h0034,-16'h0017,-16'h007e,-16'h00dc,16'h0016,16'h0182,16'h00ae,-16'h006c,16'h0015,-16'h00ce,-16'h0053,16'h0042,16'h0107,-16'h0136,16'h0058,-16'h002d,16'h0064,16'h0099,16'h00b5,-16'h00ce,-16'h0061,-16'h000b,16'h0080,-16'h0009,-16'h002f,-16'h001a,-16'h0025,-16'h0086,16'h02de,16'h009b,-16'h0095,16'h01ee,16'h001c,-16'h006f,16'h00e4,16'h004a,-16'h03e7,-16'h0292,-16'h000d,-16'h0281,-16'h0160,16'h0009,-16'h000a,-16'h0087,16'h0004,16'h00db,-16'h002c,-16'h013e,-16'h0072,16'h00bf,16'h0041,-16'h0038,-16'h002d,-16'h00b9,16'h0021,16'h003b,16'h009e,-16'h0158,16'h01fa,-16'h0019,16'h0070,-16'h0039,16'h0048,16'h0201,16'h0036,16'h0063,16'h00cf,-16'h0143,16'h0083,16'h019b,16'h00e5,16'h0042,-16'h0009,-16'h0004,-16'h0044,16'h0083,16'h00c8,16'h000d,16'h011d,-16'h0045,16'h00a9,16'h007f,16'h000a,-16'h0037,-16'h00bb,16'h0027,16'h00a4,16'h000e,-16'h0002,16'h0078,-16'h00c1,-16'h0032,16'h02c9,16'h011d,-16'h0088,16'h0220,16'h00ec,-16'h0105,16'h0160,-16'h0024,-16'h0371,-16'h0275,16'h007f,-16'h02ca,-16'h0214,-16'h000d,-16'h0040,-16'h0057,16'h0005,16'h00a2,-16'h003d,-16'h00c0,16'h0086,16'h00ba,16'h0028,-16'h0092,16'h005a,-16'h00c8,-16'h0081,16'h003f,16'h0061,-16'h00bf,16'h01a9,-16'h0065,-16'h000d,-16'h002b,16'h000a,16'h01f9,16'h0070,16'h0067,16'h020a,-16'h00e6,-16'h0021,16'h010c,16'h0110,16'h001b,-16'h0016,-16'h000f,-16'h002b,16'h0061,16'h0043,16'h00a4,16'h00e9,-16'h002a,16'h007f,16'h0017,16'h0042,16'h0028,-16'h009d,16'h000f,16'h0099,16'h003a,-16'h0037,16'h000d,-16'h0077,16'h005e,16'h0232,16'h00f3,-16'h0106,16'h0268,16'h0086,-16'h00b2,16'h008f,-16'h005f,-16'h0383,-16'h0308,16'h0023,-16'h027d,-16'h016b,16'h008f,16'h0008,16'h0000,16'h003b,16'h00d9,16'h003e,-16'h0030,16'h0055,-16'h000f,16'h0019,-16'h0053,16'h001d,-16'h007d,-16'h0073,16'h0002,16'h009d,16'h000e,16'h01d7,-16'h0066,-16'h00dc,16'h000d,16'h0040,16'h020e,16'h0051,16'h000c,16'h0174,-16'h0083,-16'h0036,-16'h008c,16'h014c,16'h0049,-16'h0024,-16'h0070,16'h003a,16'h006c,-16'h0064,16'h0138,16'h0103,-16'h005c,-16'h0043,16'h00be,16'h000f,16'h005f,-16'h0149,16'h0087,16'h00d5,-16'h003e,-16'h0097,16'h005f,-16'h0003,16'h00b4,16'h01d8,16'h011d,-16'h00d2,16'h0244,16'h00c5,-16'h010a,-16'h0008,-16'h00f2,-16'h0268,-16'h033c,16'h009f,-16'h025c,-16'h018b,16'h0024,16'h0015,-16'h0035,16'h00bf,16'h0113,16'h0068,-16'h0063,16'h00f5,-16'h0066,16'h0033,-16'h00f2,16'h0047,-16'h0066,-16'h008a,16'h0009,16'h007d,16'h002a,16'h017c,-16'h0070,-16'h0153,16'h001f,16'h0050,16'h0147,16'h004f,16'h0024,16'h0164,-16'h005a,-16'h008a,-16'h01a0,16'h00fa,16'h00d4,-16'h004b,16'h0003,16'h0033,16'h007a,-16'h0212,16'h015c,16'h0098,-16'h00cb,-16'h016c,16'h0059,-16'h006c,16'h003b,-16'h00f8,16'h0042,16'h010d,16'h0067,-16'h0097,16'h0077,-16'h0004,16'h00f9,16'h01d2,16'h00df,-16'h00e7,16'h0251,16'h0032,-16'h00e4,-16'h0067,-16'h01b1,-16'h0192,-16'h026e,16'h0075,-16'h025f,-16'h0193,-16'h0052,-16'h0027,-16'h0018,16'h0032,16'h011f,16'h0047,16'h00cd,16'h0097,-16'h006f,16'h002f,-16'h00c3,16'h007a,-16'h0002,-16'h0012,16'h0013,16'h001c,16'h0086,16'h01a1,-16'h0048,-16'h0111,-16'h003b,-16'h001e,16'h0105,-16'h008e,16'h0019,16'h00e4,16'h0096,-16'h004d,-16'h0099,16'h008d,16'h0032,-16'h00c5,16'h008b,16'h0054,16'h007e,-16'h04d7,16'h0165,16'h003c,-16'h008d,-16'h0119,16'h0024,-16'h00f9,-16'h0059,-16'h004d,16'h00a1,16'h0028,16'h001f,-16'h00c4,16'h00b2,-16'h0065,16'h0118,16'h019d,-16'h0019,-16'h0074,16'h01c6,16'h0047,-16'h0073,-16'h009a,-16'h02e7,-16'h0115,-16'h02c6,16'h00f9,-16'h026f,-16'h0191,16'h0039,16'h0040,16'h0036,16'h000b,16'h0147,16'h0056,16'h018e,16'h00fc,-16'h00e9,16'h00de,-16'h0093,16'h005a,-16'h000f,16'h0030,16'h0070,16'h0094,16'h0116,16'h01ec,-16'h001d,-16'h003c,-16'h00d9,16'h0047,16'h0010,-16'h0076,-16'h0030,16'h00de,16'h011b,-16'h00a6,-16'h003d,-16'h001b,16'h00d3,-16'h015b,-16'h0007,16'h008b,16'h0072,-16'h065d,16'h0193,16'h00a6,-16'h0047,-16'h009e,16'h0022,-16'h0019,16'h001b,16'h00e3,16'h0033,-16'h005d,16'h0028,-16'h0119,16'h0097,-16'h012d,16'h00fd,16'h018d,-16'h01e8,-16'h010e,16'h0216,16'h0020,16'h0080,-16'h0067,-16'h0375,16'h0033,-16'h022b,16'h004c,-16'h0321,-16'h0174,16'h003c,16'h005f,16'h001c,16'h0079,16'h0112,16'h00a8,16'h0191,16'h00d1,-16'h00ae,16'h00e6,-16'h0057,-16'h001e,-16'h0004,16'h0135,16'h0046,16'h0147,16'h00c5,16'h01b7,-16'h000d,16'h001c,-16'h008e,16'h001d,-16'h009a,-16'h0037,-16'h0032,16'h0092,16'h01b0,-16'h008a,16'h001d,-16'h0166,16'h00b3,-16'h014b,16'h005a,16'h007c,16'h0058,-16'h04e9,16'h0198,16'h0073,16'h0010,16'h002d,16'h006b,16'h002a,-16'h006d,16'h014d,-16'h0035,-16'h01fa,-16'h0037,-16'h00c5,16'h006d,-16'h014c,16'h006c,16'h00a5,-16'h00ff,-16'h0098,16'h0256,16'h000c,16'h0090,-16'h00ea,-16'h043b,16'h0145,-16'h027e,16'h0067,-16'h0275,-16'h01d5,16'h0078,16'h002d,16'h0032,16'h0031,16'h0095,16'h00ee,16'h0148,16'h012d,-16'h00c0,16'h0138,16'h0041,-16'h0010,16'h000b,16'h0101,16'h002a,16'h018a,16'h008c,16'h0140,16'h005b,-16'h00b3,-16'h0064,-16'h0062,-16'h01dc,16'h008b,-16'h001d,16'h0033,16'h0180,-16'h000f,-16'h005c,-16'h047a,16'h00bf,-16'h00fe,16'h0038,16'h006a,16'h006f,-16'h0249,16'h00d6,16'h00b7,16'h00d0,-16'h0039,16'h0065,16'h006d,-16'h0027,16'h00b9,-16'h0014,-16'h0294,-16'h0026,-16'h0145,16'h004f,-16'h00de,-16'h00c7,16'h0059,16'h0035,-16'h0071,16'h0223,16'h001f,16'h0124,-16'h00da,-16'h03d2,16'h017c,-16'h021f,16'h0029,-16'h0200,-16'h01a1,16'h0052,16'h0030,16'h004e,16'h0052,16'h0079,16'h0052,16'h00cd,16'h0175,-16'h0022,16'h00ed,16'h00c0,16'h0073,-16'h0012,16'h01c5,16'h002a,16'h01a1,16'h007e,16'h00dd,16'h002d,16'h0000,16'h004c,16'h0047,-16'h021a,16'h0094,-16'h0025,-16'h007e,16'h01b1,16'h00a9,-16'h0050,-16'h0514,16'h012f,-16'h000c,16'h0040,16'h001c,16'h017d,-16'h017a,16'h00ec,16'h00a1,16'h007d,16'h0042,16'h0055,16'h00cc,-16'h000c,16'h0052,-16'h00af,-16'h0246,-16'h0040,-16'h0105,-16'h0048,-16'h0076,-16'h0144,16'h0106,16'h0143,-16'h007f,16'h02a0,16'h005d,16'h00b0,-16'h0092,-16'h031a,16'h01b7,-16'h011f,-16'h0120,-16'h01a4,-16'h007f,16'h00a5,-16'h003a,16'h007a,16'h00a5,-16'h0026,16'h003b,16'h0048,16'h01b3,16'h0043,16'h0195,16'h015f,16'h0018,-16'h00a0,16'h014c,-16'h0007,16'h017f,16'h007a,16'h00ff,16'h0077,-16'h0008,16'h0034,16'h0052,-16'h0190,16'h006d,16'h008b,-16'h0205,16'h0111,16'h0110,-16'h007e,-16'h038b,16'h0119,16'h0065,16'h0039,-16'h003d,16'h00bd,-16'h0130,16'h00bd,16'h00d5,-16'h0011,-16'h00db,-16'h0070,16'h0132,-16'h002e,-16'h0077,-16'h0066,-16'h0282,-16'h0033,-16'h00fd,16'h0035,-16'h0007,-16'h0100,16'h00b9,16'h027a,-16'h00e8,16'h0267,16'h014b,16'h00ae,-16'h007b,-16'h01f8,16'h0206,-16'h0019,-16'h0118,-16'h01fa,16'h000a,16'h0105,-16'h008c,16'h0094,16'h007d,-16'h0064,16'h0064,-16'h0036,16'h015d,16'h012a,16'h016b,16'h014b,-16'h0016,-16'h00d4,16'h00f9,16'h002c,16'h016e,16'h007f,16'h0065,16'h011a,-16'h00ab,16'h006e,-16'h0032,-16'h0183,16'h009d,16'h0073,-16'h02d0,16'h00a0,16'h00b0,-16'h005d,-16'h012f,16'h0175,16'h00f6,-16'h001d,-16'h007f,16'h0044,-16'h0034,16'h0049,16'h0012,-16'h00e1,-16'h005f,-16'h005d,16'h00da,-16'h001d,-16'h00b9,-16'h00cc,-16'h014a,-16'h0022,-16'h015d,-16'h0048,16'h005c,-16'h00b9,16'h0128,16'h025f,-16'h0094,16'h0243,16'h00e9,16'h0095,-16'h0082,-16'h0111,16'h01af,16'h00f9,-16'h00e5,-16'h01f2,-16'h0039,16'h016c,-16'h003b,16'h0038,16'h005f,-16'h0181,16'h00d4,-16'h000a,16'h00e1,16'h0157,16'h0159,16'h01f0,-16'h0007,-16'h007f,16'h009f,16'h0093,16'h0151,16'h00d8,16'h005c,16'h00c4,-16'h000a,16'h0057,-16'h003b,-16'h0174,16'h0095,16'h00d5,-16'h03d9,16'h00cc,16'h0081,-16'h0079,16'h00bb,16'h016b,16'h00d1,16'h001f,-16'h00b9,16'h009b,-16'h0063,16'h002f,16'h002f,-16'h0142,-16'h010b,16'h0021,16'h009c,16'h003b,-16'h00f8,16'h00b0,-16'h00bd,-16'h0097,-16'h0188,-16'h0039,-16'h002e,-16'h0086,16'h0191,16'h01dc,-16'h005b,16'h0235,16'h0106,16'h0078,16'h0035,-16'h00c4,16'h0161,16'h014d,-16'h0092,-16'h01be,16'h000b,16'h0145,-16'h0064,-16'h003e,-16'h0036,-16'h0106,16'h00da,16'h0079,16'h002f,16'h00d7,16'h0025,16'h0174,16'h00bf,-16'h0090,16'h0094,16'h00fb,16'h00c8,16'h0093,16'h0087,16'h00a1,-16'h001d,16'h00a1,16'h001b,-16'h00eb,16'h00bb,16'h00fd,-16'h0371,16'h00ea,16'h0101,-16'h008e,16'h00c7,16'h0105,16'h0126,-16'h008a,-16'h0064,16'h003e,-16'h002a,16'h0001,-16'h0004,-16'h015c,-16'h0115,16'h0013,16'h0024,-16'h0075,-16'h00f6,16'h0108,-16'h00ab,-16'h007e,-16'h01bf,-16'h002a,-16'h003d,-16'h0065,16'h026c,16'h00ec,16'h0024,16'h018f,16'h013c,16'h00c3,16'h00c8,-16'h0041,16'h0175,16'h0101,16'h000c,-16'h018d,16'h0009,16'h014d,-16'h002f,-16'h003b,-16'h0009,-16'h00d6,16'h0062,16'h0013,16'h0032,16'h00d4,-16'h0073,16'h015c,16'h00a0,-16'h0063,16'h0054,16'h00a5,16'h00d0,16'h00c0,16'h00bf,16'h006a,-16'h0034,16'h00ac,-16'h0031,-16'h011d,16'h0065,16'h0062,-16'h02d9,16'h0025,16'h00c3,16'h0030,16'h00fc,16'h0132,16'h00d7,16'h0043,16'h0018,16'h00be,16'h0040,-16'h0006,-16'h0066,-16'h00f9,-16'h012a,16'h00c9,16'h004a,16'h001c,-16'h00c9,16'h009c,-16'h006d,-16'h0069,-16'h014f,-16'h0027,16'h0029,-16'h0062,16'h023e,16'h006c,16'h0018,16'h00ab,16'h01b5,16'h0055,16'h0105,-16'h006f,16'h016f,16'h0112,16'h0033,-16'h0138,16'h00c2,16'h01b6,-16'h0106,16'h0012,16'h0078,-16'h0088,16'h006e,-16'h000d,16'h003c,16'h0019,-16'h0131,16'h01b5,16'h00fd,-16'h0016,16'h0015,-16'h003d,-16'h00b3,-16'h00cc,16'h00ef,16'h0015,-16'h0080,16'h0038,16'h022a,-16'h01ad,16'h00be,16'h0080,16'h004a,16'h0042,-16'h0096,-16'h01de,16'h00fe,16'h0219,-16'h0009,16'h000e,-16'h0006,16'h00b8,-16'h0087,-16'h000f,16'h01bf,16'h00de,-16'h00a8,16'h0163,16'h003f,16'h0017,16'h001d,-16'h0022,-16'h0177,-16'h00f5,-16'h0072,-16'h0012,-16'h0046,16'h005e,16'h0129,16'h00a9,16'h0006,16'h00fb,-16'h00b7,16'h01d8,16'h0016,16'h0103,-16'h004d,-16'h0100,16'h00e9,-16'h00a2,16'h00a6,-16'h0163,-16'h0071,-16'h010e,-16'h00a8,16'h0009,16'h016f,-16'h00fd,16'h00a9,-16'h00d1,16'h0080,-16'h008a,-16'h0028,-16'h00fe,-16'h00a1,16'h0001,-16'h00f5,-16'h00ae,16'h0138,-16'h0059,-16'h005e,16'h0048,16'h0208,-16'h02da,16'h0179,16'h0068,16'h000e,16'h00d9,-16'h0031,-16'h0178,16'h00d9,16'h015d,16'h006e,16'h0044,-16'h0036,16'h00c5,-16'h00e4,-16'h00ea,16'h02c1,16'h0091,-16'h00ad,16'h00d5,16'h0023,-16'h0008,16'h006a,16'h003e,-16'h00e8,-16'h00cc,-16'h0012,16'h0021,-16'h0052,16'h0033,16'h0205,16'h0166,16'h0040,16'h00b0,-16'h008a,16'h01c1,16'h0145,16'h00e7,-16'h00a3,-16'h001e,16'h0067,-16'h0035,16'h00ea,-16'h01bd,-16'h017d,-16'h00b1,-16'h009c,-16'h0083,16'h0144,-16'h0096,16'h0154,-16'h0066,16'h0006,-16'h0042,-16'h0014,-16'h016a,-16'h00c4,16'h0034,-16'h01af,-16'h0073,16'h0185,-16'h005c,-16'h00c0,-16'h0036,16'h00fa,-16'h02b5,16'h00fe,16'h00b9,-16'h00be,16'h0186,-16'h0014,-16'h0125,16'h00bd,16'h00d4,16'h010d,16'h0029,-16'h00bb,16'h0115,-16'h012a,-16'h00ec,16'h02fb,16'h00ac,-16'h0032,16'h00c3,-16'h0006,-16'h0069,16'h002c,16'h0060,-16'h00b4,-16'h003e,-16'h0026,16'h0026,-16'h010a,16'h0077,16'h01bb,16'h0063,-16'h0048,16'h00b6,-16'h0176,16'h018a,16'h00d3,16'h0075,-16'h00c4,-16'h0015,16'h0102,-16'h0081,16'h00a5,-16'h02d7,-16'h0217,-16'h0112,-16'h0068,-16'h0080,16'h0121,-16'h00ae,16'h0140,-16'h0013,16'h001c,16'h0002,-16'h0002,-16'h00f8,-16'h0021,16'h00ed,-16'h0265,-16'h00cd,16'h026e,-16'h00c8,-16'h0105,16'h0076,16'h00e6,-16'h020f,16'h004f,16'h0147,-16'h021c,16'h013b,16'h003e,16'h0046,16'h00c2,16'h0012,16'h0083,16'h0021,-16'h00da,16'h0101,-16'h00bf,-16'h0131,16'h018f,16'h0091,-16'h009d,16'h0141,-16'h0071,16'h001f,-16'h008f,16'h002f,16'h000b,-16'h0077,-16'h008e,16'h0055,-16'h0128,-16'h0046,16'h020b,-16'h000e,16'h009d,16'h00de,-16'h011b,16'h00ab,16'h008a,16'h00a6,-16'h00dd,16'h0010,16'h006a,-16'h005e,16'h0167,-16'h030c,-16'h028d,-16'h012f,16'h0022,-16'h00c6,16'h01ae,16'h0011,16'h0155,16'h00cc,16'h005e,16'h0022,-16'h00a3,-16'h00cc,-16'h00dc,16'h0172,-16'h0345,-16'h0053,16'h028a,-16'h0130,-16'h0090,16'h00ce,16'h005c,-16'h019b,16'h004d,16'h0055,-16'h0337,16'h01fb,16'h006f,16'h0120,16'h00d0,-16'h0094,16'h00b0,-16'h000b,-16'h00a4,16'h00a9,-16'h0019,-16'h0102,16'h0069,16'h005f,-16'h0078,16'h0143,-16'h008c,16'h0071,-16'h0045,16'h001a,16'h0048,16'h0011,-16'h0117,16'h0078,-16'h0135,16'h0060,16'h029e,16'h0028,16'h016e,16'h0102,16'h0004,16'h007b,16'h0063,16'h00cf,-16'h00f1,16'h0057,16'h0057,-16'h0148,16'h01f2,-16'h0299,-16'h01d4,-16'h0129,16'h007a,-16'h004b,16'h019e,16'h002f,16'h0164,16'h00f1,16'h0032,-16'h0001,16'h000f,-16'h006c,-16'h0088,16'h01b0,-16'h0333,16'h00a6,16'h0202,-16'h00e4,-16'h0052,16'h00f3,16'h0056,-16'h004d,16'h0010,-16'h009d,-16'h02dc,16'h01cc,16'h003a,16'h00aa,16'h0031,-16'h017e,16'h00fa,-16'h0059,-16'h00b9,16'h012e,16'h0074,-16'h011d,-16'h017e,-16'h0002,-16'h0089,16'h015f,-16'h00ec,16'h0012,-16'h0043,-16'h001e,16'h013d,-16'h001c,-16'h00d9,-16'h003f,-16'h00b8,16'h007f,16'h02e9,-16'h003b,16'h016c,16'h011f,16'h005e,16'h009e,16'h0035,16'h00c4,-16'h0130,-16'h00a0,16'h006d,-16'h0216,16'h01d2,-16'h023b,-16'h003d,-16'h00f6,16'h00bb,-16'h0078,16'h01e5,16'h015f,16'h0111,16'h013a,-16'h001b,16'h0013,16'h0024,-16'h004f,-16'h0030,16'h01ba,-16'h01d2,16'h0102,16'h0251,-16'h007e,-16'h0091,16'h0093,-16'h005f,-16'h002b,-16'h004a,-16'h00d9,-16'h0327,16'h01e0,16'h0041,16'h0016,16'h0016,-16'h0142,16'h013b,-16'h006c,-16'h003b,16'h00dc,16'h0007,-16'h018b,-16'h039e,16'h0096,16'h003d,16'h011e,-16'h0049,-16'h0025,16'h000c,16'h003c,16'h0107,-16'h00d0,-16'h0159,16'h0001,16'h0086,16'h0074,16'h029b,-16'h0037,16'h0146,16'h012c,16'h00f7,16'h0097,16'h00f2,16'h004f,-16'h019b,-16'h0040,16'h0052,-16'h0290,16'h011a,-16'h014c,-16'h0073,-16'h0145,16'h013a,-16'h0042,16'h011c,16'h011a,16'h011b,16'h012c,16'h002a,-16'h0063,16'h003c,-16'h0034,-16'h003c,16'h01a0,-16'h0072,16'h00df,16'h0282,-16'h006b,-16'h006c,16'h005b,-16'h0027,16'h0045,-16'h0065,-16'h009d,-16'h01f2,16'h0109,-16'h002f,-16'h0081,-16'h0026,-16'h00b0,16'h00cc,-16'h0063,-16'h004b,16'h001a,16'h000c,-16'h016c,-16'h04a8,16'h010c,-16'h0002,16'h0116,-16'h0090,-16'h0016,-16'h00b8,16'h000b,16'h0190,-16'h0054,-16'h010e,-16'h006b,16'h0162,-16'h0017,16'h025d,-16'h00a1,16'h0169,16'h0141,16'h00a6,16'h0132,16'h012e,16'h0017,-16'h013b,16'h002d,-16'h0087,-16'h02ab,16'h0072,16'h0030,16'h000e,-16'h012e,16'h00ab,-16'h005c,16'h0084,16'h0160,16'h0134,16'h0133,-16'h004a,-16'h0038,-16'h000a,-16'h0078,-16'h0089,16'h01bd,16'h0000,16'h0096,16'h027c,-16'h007c,-16'h00c1,16'h0042,-16'h00b0,16'h0046,-16'h006e,-16'h0068,-16'h0230,16'h00fe,-16'h003b,-16'h0106,16'h0068,-16'h0164,16'h0111,-16'h0009,16'h003e,16'h00bd,16'h002d,-16'h0224,-16'h04cb,16'h00bb,16'h0024,16'h006a,-16'h0091,-16'h0066,-16'h0060,-16'h0042,16'h017c,-16'h0001,-16'h003d,-16'h001c,16'h00de,-16'h00be,16'h02af,-16'h0106,16'h0179,16'h00d9,16'h0088,16'h008d,16'h00af,16'h003e,-16'h025a,16'h0040,-16'h0071,-16'h0280,-16'h0105,16'h0059,-16'h0023,-16'h01b0,16'h007c,-16'h003a,-16'h0008,16'h0153,16'h0113,16'h00dd,-16'h007c,16'h0001,16'h007f,-16'h0091,-16'h00ba,16'h00f3,16'h0082,16'h0034,16'h0255,-16'h009b,16'h0000,-16'h002c,-16'h005f,16'h0121,-16'h0026,-16'h00ec,-16'h0199,16'h0012,-16'h0018,-16'h00f8,16'h000f,-16'h0173,16'h007a,-16'h0047,-16'h0005,16'h0044,16'h0099,-16'h01db,-16'h032c,16'h0010,-16'h004a,16'h0040,-16'h0085,16'h000c,-16'h0084,-16'h0067,16'h015d,-16'h00a7,-16'h008c,16'h002e,16'h01b4,-16'h000c,16'h02fa,-16'h004e,16'h0100,16'h0127,16'h0077,16'h00b5,16'h0113,-16'h0051,-16'h03ad,16'h0044,-16'h0044,-16'h02db,-16'h0100,16'h00ac,-16'h0057,-16'h01d7,16'h003c,-16'h0069,16'h0032,-16'h000b,16'h0049,16'h013c,-16'h0077,-16'h0061,-16'h0024,-16'h0079,-16'h00aa,16'h000f,16'h012d,-16'h0098,16'h01c2,-16'h008c,16'h0082,-16'h0068,16'h002b,16'h01ad,16'h006f,-16'h00dd,-16'h0130,-16'h00b5,-16'h0062,-16'h002c,16'h004e,-16'h0102,16'h0001,-16'h0080,16'h002d,16'h0060,16'h010a,-16'h01a4,-16'h0150,16'h0057,16'h002d,16'h004f,16'h004d,-16'h007d,-16'h003f,-16'h0055,16'h01a3,-16'h0062,16'h004d,16'h0081,16'h01eb,16'h0054,16'h024b,-16'h0021,16'h00d0,16'h0102,16'h0014,16'h00b9,16'h0144,16'h0006,-16'h057b,16'h002e,-16'h0003,-16'h0383,-16'h0042,16'h0045,-16'h0002,-16'h01b9,16'h0052,-16'h0064,16'h001e,-16'h0105,16'h0067,16'h00da,-16'h0092,-16'h0078,16'h0032,-16'h0046,16'h000c,-16'h0014,16'h00cc,-16'h00e7,16'h016e,16'h0004,16'h0084,-16'h0069,-16'h000c,16'h01b7,16'h0066,-16'h00b0,-16'h00e9,-16'h008d,-16'h0044,16'h0074,-16'h0051,-16'h00d8,-16'h0032,-16'h0011,16'h000f,16'h007a,16'h0168,-16'h0137,-16'h0012,16'h00bd,-16'h001a,16'h005c,16'h0009,-16'h0049,16'h0086,-16'h0091,16'h00c1,-16'h0002,-16'h0029,16'h00ab,16'h00a2,16'h0060,16'h0254,-16'h0053,16'h00f7,16'h0126,16'h0049,16'h0077,16'h00c0,-16'h0004,-16'h0511,-16'h0047,-16'h0018,-16'h030e,-16'h0099,-16'h004a,-16'h004c,-16'h0147,16'h0002,16'h0063,16'h0044,-16'h0168,16'h0090,16'h007f,16'h0008,-16'h0095,-16'h0010,-16'h006b,16'h005b,-16'h0097,16'h00f7,-16'h009d,16'h01dc,16'h0031,16'h00b9,-16'h0045,16'h002f,16'h01dc,-16'h0014,-16'h0009,-16'h00f3,-16'h0157,-16'h0037,16'h0162,16'h005a,-16'h00d9,-16'h000f,-16'h004d,-16'h0036,16'h00d4,16'h0161,-16'h0122,16'h00fd,-16'h000b,-16'h0031,16'h0047,16'h005a,-16'h0018,16'h007e,-16'h006b,16'h00fb,-16'h0035,-16'h0062,16'h0041,-16'h003d,-16'h0047,16'h0272,16'h001a,16'h00ac,16'h0187,16'h0096,-16'h0055,16'h018f,16'h0006,-16'h0352,-16'h0069,16'h0050,-16'h0341,-16'h00d0,-16'h0005,-16'h0020,-16'h0140,-16'h0054,16'h00b4,16'h0000,-16'h016d,16'h0028,16'h0092,16'h0015,-16'h0097,-16'h0046,-16'h00a2,16'h003b,-16'h00bd,16'h0092,-16'h006f,16'h021a,16'h0034,16'h00c3,-16'h0070,16'h0001,16'h0215,-16'h0025,-16'h0070,-16'h0064,-16'h0101,16'h0032,16'h0185,16'h00c8,-16'h006d,-16'h0006,-16'h00a6,-16'h0014,16'h00b5,16'h0119,-16'h000a,16'h016a,-16'h0005,16'h0018,16'h0061,16'h0031,-16'h0078,16'h0024,-16'h0054,16'h00b7,-16'h003f,-16'h00cc,-16'h0011,-16'h0073,-16'h00a2,16'h02a3,16'h008c,16'h00af,16'h026c,16'h007a,16'h000d,16'h00e2,-16'h002a,-16'h0214,-16'h0102,16'h0062,-16'h034f,-16'h015b,-16'h0028,-16'h0067,-16'h0196,-16'h0080,16'h00e7,16'h0032,-16'h00b0,16'h00c5,16'h0032,16'h0051,-16'h008a,16'h0011,-16'h0028,16'h00a2,16'h0000,16'h0043,-16'h0066,16'h0205,16'h003b,16'h0053,-16'h0001,16'h0034,16'h023c,16'h0036,16'h0030,16'h006f,-16'h00d9,16'h0010,16'h0140,16'h0120,-16'h001b,16'h006f,-16'h0027,-16'h0031,16'h0093,16'h0146,16'h00b6,16'h0149,16'h0063,16'h0034,16'h0039,-16'h0015,-16'h0023,16'h0038,-16'h0025,16'h00b1,-16'h008e,-16'h006c,-16'h0060,-16'h014b,-16'h0092,16'h028b,16'h008d,16'h00e3,16'h0295,16'h00ae,-16'h00ed,16'h0138,-16'h0057,-16'h0244,-16'h00d2,16'h0087,-16'h030f,-16'h01f8,16'h0043,-16'h004b,-16'h01e5,16'h0036,16'h008b,-16'h0068,-16'h0078,16'h00a7,-16'h0027,-16'h0046,-16'h00b7,16'h002b,-16'h00bf,-16'h0042,16'h0003,16'h00d2,16'h0031,16'h0259,-16'h004d,-16'h003d,-16'h0048,16'h0027,16'h0208,16'h006e,16'h005d,16'h0198,-16'h00ce,16'h0032,-16'h004d,16'h00f9,16'h0018,16'h00ea,-16'h0077,-16'h0071,16'h00cd,16'h009c,16'h0129,16'h01bd,-16'h0036,16'h0002,16'h0003,16'h002c,16'h0046,-16'h00bb,-16'h0038,16'h008b,-16'h0049,-16'h007b,16'h0089,-16'h0083,-16'h0029,16'h021e,16'h00c1,16'h00cd,16'h028c,16'h003d,-16'h00b1,16'h00e8,16'h008f,-16'h0234,-16'h01db,16'h011c,-16'h0307,-16'h0171,16'h00bd,-16'h008b,-16'h0136,16'h0034,16'h0100,-16'h0013,16'h00ac,16'h009f,-16'h0006,-16'h000e,-16'h00ef,16'h0051,-16'h007c,-16'h00c8,16'h003e,16'h00b0,16'h0042,16'h0210,-16'h0085,16'h0006,-16'h003a,16'h0052,16'h0177,16'h002b,16'h0014,16'h0185,-16'h0088,-16'h0018,-16'h021b,16'h01b8,16'h00b2,16'h0085,-16'h0024,16'h0035,16'h0098,-16'h0090,16'h018b,16'h0141,16'h0056,-16'h008a,16'h0077,16'h0019,16'h0026,-16'h00f1,-16'h001c,16'h00af,16'h0047,-16'h0083,16'h003e,-16'h0054,16'h0081,16'h0231,16'h012e,16'h009c,16'h02c2,16'h000c,-16'h00f2,16'h0049,-16'h0031,-16'h017d,-16'h01ec,16'h0105,-16'h035f,-16'h017b,16'h0081,-16'h006e,-16'h0167,16'h0035,16'h015f,16'h0032,16'h00cb,16'h00e7,-16'h0096,16'h0010,-16'h00e3,16'h004a,-16'h0007,-16'h0058,-16'h000c,16'h011f,16'h007c,16'h0141,-16'h00a0,-16'h0077,-16'h0027,-16'h0001,16'h0059,-16'h000f,16'h0064,16'h017c,-16'h00a5,-16'h0051,-16'h01d4,16'h010e,16'h0110,-16'h003e,16'h003a,-16'h0015,16'h00a7,-16'h0207,16'h0193,16'h0088,-16'h004e,-16'h0128,16'h0024,-16'h003b,16'h001b,-16'h0148,-16'h0004,16'h0040,16'h00b6,-16'h0039,16'h00bf,16'h0011,16'h00e2,16'h022a,16'h010d,16'h0057,16'h024e,16'h0062,-16'h011c,-16'h0090,-16'h0179,-16'h00c2,-16'h0250,16'h00ca,-16'h0344,-16'h0111,16'h001c,-16'h0016,-16'h00fb,16'h00c6,16'h0185,16'h0040,16'h0118,16'h012a,-16'h0118,16'h0096,-16'h00d2,16'h000c,-16'h005e,16'h0009,-16'h000a,16'h0111,16'h011e,16'h0153,-16'h0098,-16'h0059,-16'h010a,16'h004f,-16'h002c,-16'h0055,16'h0031,16'h019e,16'h0099,-16'h0043,-16'h012e,16'h0149,16'h01b7,-16'h0041,16'h0046,16'h004b,16'h0122,-16'h0569,16'h01ca,16'h002e,-16'h000f,-16'h0108,-16'h0079,-16'h0027,-16'h009b,-16'h0074,-16'h0035,-16'h004a,16'h00b8,16'h0004,16'h00b6,-16'h0089,16'h0159,16'h0207,-16'h0041,16'h0080,16'h0199,-16'h005e,-16'h0085,-16'h0068,-16'h026f,16'h002e,-16'h0268,16'h0125,-16'h02b8,-16'h0145,16'h0045,-16'h0077,-16'h00ea,16'h0060,16'h0196,16'h004f,16'h013e,16'h0103,-16'h00d5,16'h00c8,-16'h0049,16'h0009,16'h004b,16'h00b2,16'h0054,16'h0104,16'h011a,16'h01bc,-16'h00c6,-16'h000d,-16'h0171,-16'h0063,-16'h00b2,-16'h0085,16'h0061,16'h01b8,16'h00ea,-16'h003c,-16'h00a6,16'h0026,16'h01b6,-16'h014e,16'h0023,-16'h0008,16'h011a,-16'h07be,16'h013e,16'h0041,-16'h000f,-16'h00ad,16'h0041,16'h002a,-16'h0088,16'h0014,-16'h0003,-16'h0102,-16'h0002,16'h0047,16'h00ed,-16'h0140,16'h0111,16'h01af,-16'h0254,16'h0023,16'h0200,-16'h0001,-16'h0025,-16'h00b2,-16'h03f9,16'h013e,-16'h0233,16'h00df,-16'h0305,-16'h01dd,16'h0058,-16'h003a,-16'h0096,16'h0078,16'h0166,16'h00f8,16'h00ee,16'h00cb,-16'h0028,16'h00d7,-16'h002d,16'h0012,16'h0000,16'h016b,-16'h0057,16'h01df,16'h0135,16'h00dc,-16'h001a,16'h004a,-16'h00db,-16'h0010,-16'h018a,16'h002d,16'h0063,16'h0103,16'h014b,16'h008e,16'h0037,-16'h011e,16'h0194,-16'h01c6,16'h0026,16'h009b,16'h0084,-16'h0545,16'h0129,16'h0039,-16'h0073,-16'h004f,-16'h0004,16'h007b,-16'h0071,16'h01b2,16'h0023,-16'h01d2,-16'h0037,16'h0040,16'h00af,-16'h011c,16'h00cf,16'h00ca,-16'h01e9,16'h0072,16'h01ff,16'h004d,16'h0106,-16'h00c0,-16'h04a6,16'h01f5,-16'h02e4,16'h00b6,-16'h02fc,-16'h0194,16'h0036,16'h0047,-16'h0007,16'h0082,16'h0162,16'h00e4,16'h00c6,16'h0135,16'h0030,16'h0181,16'h0023,16'h0026,16'h0022,16'h014e,-16'h00a3,16'h01e2,16'h018b,16'h0101,-16'h0040,16'h00a1,-16'h012e,16'h0016,-16'h02b2,-16'h0038,16'h0043,16'h00d3,16'h0147,16'h010c,16'h0007,-16'h033c,16'h01e3,-16'h0110,16'h004a,16'h0083,16'h00c3,-16'h0279,16'h0059,-16'h0018,16'h0107,-16'h0026,16'h008f,16'h0098,-16'h005b,16'h0178,16'h0008,-16'h0295,-16'h005b,-16'h0036,16'h009c,-16'h00e5,16'h0000,16'h0094,16'h004d,16'h0076,16'h01b9,16'h0001,16'h0195,-16'h007b,-16'h040b,16'h01df,-16'h02e1,16'h0056,-16'h0342,-16'h0035,16'h0008,16'h0062,-16'h0021,16'h003a,16'h0120,16'h00f1,16'h003e,16'h015b,16'h002a,16'h0154,16'h009c,16'h006c,-16'h0016,16'h0156,16'h002a,16'h021a,16'h00e9,16'h00f2,16'h005a,16'h0057,-16'h0039,16'h0004,-16'h02ef,16'h0076,16'h008e,16'h0028,16'h0144,16'h00e6,-16'h006f,-16'h046a,16'h014c,-16'h00c0,16'h001c,16'h006f,16'h00d4,-16'h01d6,16'h0041,16'h0087,16'h006e,-16'h003c,-16'h0027,16'h0134,-16'h009b,16'h0089,-16'h0020,-16'h02f1,16'h0006,-16'h00ec,16'h0065,-16'h0045,-16'h0104,16'h00c9,16'h0208,16'h0069,16'h01f9,16'h0089,16'h0121,-16'h0084,-16'h038f,16'h024a,-16'h01d0,-16'h002d,-16'h028d,16'h002f,16'h000f,16'h0003,-16'h0080,16'h00da,16'h00bf,16'h003c,-16'h0063,16'h0211,16'h004d,16'h017a,16'h0153,16'h0092,-16'h003f,16'h01c0,16'h0019,16'h01be,16'h009a,16'h0099,16'h00a8,16'h00b6,16'h0063,16'h007c,-16'h036d,16'h002a,16'h00b0,-16'h00ed,16'h0164,16'h0066,16'h0019,-16'h0326,16'h01cb,16'h002e,16'h006a,16'h002d,16'h0144,-16'h00b4,16'h0083,16'h0008,-16'h000f,16'h0011,-16'h0085,16'h00cd,-16'h00e5,-16'h00a6,-16'h003c,-16'h0248,-16'h0068,-16'h021c,16'h0080,-16'h0004,-16'h01ae,16'h00d9,16'h02d2,16'h0010,16'h01d4,16'h0093,16'h00bc,-16'h0059,-16'h025c,16'h01ed,-16'h0117,-16'h0062,-16'h01ec,16'h0095,16'h00c8,-16'h008d,16'h001e,16'h0069,-16'h0046,16'h003a,-16'h00ca,16'h0250,16'h00de,16'h0164,16'h022b,-16'h0056,-16'h0044,16'h0102,16'h005d,16'h0113,16'h00b9,16'h00c5,16'h0088,16'h00f0,16'h0047,-16'h005d,-16'h0267,16'h0051,16'h0173,-16'h0268,16'h0111,16'h00c1,-16'h0010,-16'h016c,16'h018f,16'h00b5,16'h006b,16'h0054,16'h0079,-16'h0066,16'h00b4,-16'h004c,-16'h004a,-16'h0080,-16'h00c9,16'h0107,-16'h0089,-16'h00d4,-16'h00b1,-16'h01b7,-16'h0050,-16'h023d,16'h008f,-16'h003b,-16'h012c,16'h0141,16'h02dd,16'h002f,16'h01c7,16'h0108,16'h011b,-16'h0087,-16'h0161,16'h0232,-16'h001e,-16'h0102,-16'h01d3,16'h00d1,16'h00f8,-16'h00f7,16'h006f,16'h002c,-16'h01df,16'h0091,-16'h00d5,16'h0180,16'h00a8,16'h014b,16'h01f9,-16'h0050,-16'h0090,16'h00c4,16'h005b,16'h0119,16'h00ce,16'h002a,16'h00e0,16'h00b7,16'h00b6,16'h0049,-16'h020d,16'h006c,16'h0166,-16'h0372,16'h00f3,16'h00ca,-16'h0032,16'h007a,16'h0119,16'h00d6,16'h0055,-16'h0040,16'h0093,-16'h0002,-16'h000b,-16'h00d9,-16'h00f3,-16'h0121,16'h0033,16'h0091,-16'h00e2,-16'h0137,-16'h0048,-16'h0120,-16'h0082,-16'h02b4,16'h0009,-16'h0073,-16'h012b,16'h01da,16'h0276,16'h0046,16'h0182,16'h0104,16'h00e2,16'h000e,-16'h0085,16'h0160,16'h0039,-16'h0070,-16'h0153,16'h00cb,16'h00c5,16'h0004,16'h0047,-16'h00b3,-16'h01a1,16'h006d,-16'h0044,16'h00f9,16'h0133,16'h00f7,16'h01fb,16'h0005,-16'h00a2,16'h0057,16'h0072,16'h0030,16'h00fd,-16'h002c,16'h00e8,16'h0043,16'h0069,-16'h002c,-16'h017d,16'h00d6,16'h00bf,-16'h043c,16'h0174,16'h00db,-16'h0013,16'h0142,16'h0114,16'h016c,-16'h005e,-16'h00c2,16'h0032,-16'h0059,-16'h006b,-16'h00ca,-16'h0127,-16'h00f8,16'h006b,16'h001e,-16'h0075,-16'h01c1,16'h00e5,-16'h00a8,16'h0034,-16'h0233,16'h002e,-16'h0013,-16'h0087,16'h020f,16'h012b,16'h00a8,16'h0154,16'h013d,16'h0133,16'h0091,-16'h005f,16'h0113,16'h0132,16'h0025,-16'h013d,16'h007b,16'h00f7,-16'h0053,16'h0039,-16'h00f4,-16'h0204,16'h0098,16'h003e,16'h0030,16'h00e0,-16'h0057,16'h0193,-16'h0011,-16'h0013,-16'h0052,16'h00ec,16'h004a,16'h00b2,16'h00ae,16'h00ab,16'h0000,16'h00a0,-16'h000a,-16'h010b,16'h00e9,16'h0093,-16'h03b8,16'h0098,16'h010e,16'h004f,16'h014b,16'h0165,16'h014b,16'h0040,-16'h0085,16'h0070,-16'h0057,-16'h004e,-16'h007f,-16'h00e8,-16'h0074,16'h004a,16'h00a6,-16'h0083,-16'h0150,16'h0190,-16'h00ba,16'h001f,-16'h01d3,16'h0024,16'h000d,-16'h0003,16'h0250,16'h0080,16'h0035,16'h00a2,16'h019d,16'h00af,16'h017a,-16'h0054,16'h008d,16'h00ec,16'h0024,-16'h00a9,16'h0116,16'h01bb,-16'h0082,16'h0003,-16'h0074,-16'h01a9,16'h005a,-16'h0058,16'h0078,16'h0067,-16'h01b1,16'h01eb,16'h003a,-16'h00a7,-16'h004d,16'h0036,-16'h00cf,-16'h016f,16'h005c,-16'h0037,-16'h00f6,16'h0074,16'h01f9,-16'h0188,16'h00b5,16'h005c,16'h0096,16'h00b0,-16'h0062,-16'h0213,16'h00f6,16'h01f7,-16'h0008,16'h006d,16'h0032,16'h00e1,-16'h00fa,-16'h0036,16'h0275,16'h008c,-16'h0054,16'h015b,16'h000f,-16'h0030,16'h0036,16'h0088,-16'h00fc,-16'h0069,-16'h0019,-16'h007c,-16'h0034,16'h005f,16'h011f,16'h010c,16'h0078,16'h00d1,-16'h0095,16'h01fc,16'h00b3,16'h00fd,-16'h0078,-16'h00bf,16'h00f0,-16'h00bd,16'h00a3,-16'h0186,-16'h00c5,-16'h00b6,-16'h00d1,16'h0056,16'h0172,-16'h0135,16'h0127,-16'h00d3,16'h0023,-16'h00df,16'h005a,-16'h00c0,-16'h00ac,16'h003a,-16'h0114,-16'h00d5,16'h014a,-16'h0081,-16'h0071,16'h003b,16'h0199,-16'h0214,16'h0103,16'h005a,-16'h008c,16'h0133,16'h00a0,-16'h021c,16'h00ad,16'h010c,16'h0119,16'h003d,-16'h0078,16'h0073,-16'h0100,-16'h00ab,16'h02df,16'h00c6,-16'h0024,16'h00ec,16'h0024,-16'h0036,16'h0067,16'h0089,-16'h0134,-16'h00c2,16'h0064,-16'h0011,-16'h010e,16'h0070,16'h00e1,16'h0099,16'h012a,16'h00bb,-16'h00c2,16'h017b,16'h005e,16'h0100,-16'h00ba,-16'h0023,16'h00f7,-16'h003d,16'h008c,-16'h028e,-16'h0165,-16'h0096,16'h000f,16'h0004,16'h0116,-16'h00a9,16'h011d,16'h0054,16'h0023,-16'h0098,16'h000f,-16'h011d,-16'h00a3,16'h0083,-16'h01a3,-16'h00c5,16'h017d,-16'h00c6,-16'h00a3,16'h0035,16'h014a,-16'h027f,16'h00d7,16'h00f4,-16'h0198,16'h00fe,16'h0027,-16'h0083,16'h0113,16'h00d1,16'h00ab,-16'h0018,-16'h00d2,16'h0137,-16'h00b8,-16'h00c8,16'h026f,16'h010e,-16'h006d,16'h016b,16'h000a,-16'h007b,-16'h00b6,16'h00de,-16'h0095,-16'h0081,-16'h0009,16'h0017,-16'h0189,-16'h0066,16'h0174,16'h00ac,16'h01b6,16'h007a,-16'h018d,16'h00c0,16'h0051,16'h014c,-16'h00c8,-16'h0024,16'h00d4,-16'h00ca,16'h017b,-16'h0293,-16'h0221,-16'h0057,-16'h0022,16'h0031,16'h0122,16'h000c,16'h010c,16'h005b,16'h002d,-16'h004e,16'h002d,-16'h00e6,-16'h0073,16'h0157,-16'h029c,-16'h007a,16'h018b,-16'h00d9,-16'h0054,16'h009b,16'h00b0,-16'h01d6,16'h005f,16'h0100,-16'h02b4,16'h0124,16'h0016,16'h00b6,16'h00d0,16'h000b,16'h010f,-16'h002d,-16'h00fa,16'h0151,-16'h00cf,-16'h00f3,16'h00b0,16'h0044,-16'h000d,16'h016a,16'h0035,-16'h0048,-16'h00b3,-16'h0022,-16'h0051,-16'h008f,-16'h003d,-16'h0026,-16'h0150,-16'h0048,16'h01cd,16'h0031,16'h01e0,16'h010b,-16'h00f1,16'h00a9,16'h008d,16'h0083,-16'h0206,-16'h002b,16'h00e6,-16'h00d1,16'h022b,-16'h0228,-16'h0164,-16'h0066,16'h0006,-16'h008f,16'h0177,16'h004b,16'h017d,16'h011d,16'h00ae,16'h0013,16'h0059,-16'h00b6,-16'h014c,16'h0140,-16'h0356,16'h0042,16'h0125,-16'h00ef,-16'h0016,16'h00ec,16'h0076,-16'h0125,-16'h0035,16'h00cd,-16'h0225,16'h0182,16'h001f,16'h0137,16'h0082,-16'h0061,16'h0105,-16'h00ab,-16'h0093,16'h010c,-16'h0093,-16'h00b7,-16'h0079,16'h0028,-16'h001e,16'h0143,-16'h003a,16'h001e,-16'h0037,16'h0026,16'h009c,-16'h0086,-16'h0004,-16'h009c,-16'h0149,16'h0062,16'h024b,16'h004e,16'h01de,16'h011d,-16'h0077,16'h00dd,16'h00aa,16'h008a,-16'h0180,16'h0039,16'h005a,-16'h01dd,16'h0222,-16'h019f,-16'h00e1,16'h0010,16'h008d,-16'h0062,16'h010d,16'h00e7,16'h0137,16'h0155,-16'h0030,-16'h0019,16'h004e,-16'h00c2,-16'h0052,16'h01b6,-16'h02bd,16'h00c9,16'h01bb,-16'h00b8,-16'h0015,16'h015a,16'h0047,-16'h003f,16'h0030,16'h0001,-16'h02a1,16'h01a2,-16'h001f,16'h0044,16'h005a,-16'h0052,16'h0139,-16'h0011,-16'h007a,16'h014c,16'h0037,-16'h0115,-16'h0266,16'h0050,-16'h0003,16'h0150,-16'h0065,-16'h000c,-16'h0056,16'h0016,16'h0149,-16'h0023,16'h0020,-16'h009c,-16'h0033,16'h003c,16'h0276,-16'h003c,16'h0289,16'h0122,16'h010a,16'h00fc,16'h00c6,16'h00ea,-16'h01fb,16'h007c,-16'h0029,-16'h026d,16'h01b4,-16'h00d4,16'h0007,16'h00ab,16'h005e,-16'h00c0,16'h00bc,16'h00bf,16'h00e1,16'h00a5,-16'h0011,-16'h0014,16'h005d,-16'h001a,-16'h0036,16'h020a,-16'h0187,16'h00f4,16'h017a,-16'h0084,-16'h007a,16'h006d,-16'h0020,16'h0018,16'h004b,16'h0034,-16'h01f6,16'h014a,-16'h0066,-16'h0018,16'h0049,-16'h00d0,16'h0196,-16'h0059,-16'h0031,16'h00a9,-16'h0049,-16'h00bd,-16'h0402,16'h0121,16'h0063,16'h0113,-16'h0054,16'h0016,-16'h004f,-16'h001c,16'h01ad,-16'h001a,-16'h002d,-16'h0099,16'h00d6,-16'h0009,16'h02bb,16'h0015,16'h0293,16'h00aa,16'h00ba,16'h00e3,16'h00cb,16'h0076,-16'h01a0,16'h0075,-16'h00db,-16'h0333,16'h00af,-16'h0065,16'h000f,16'h0099,16'h009e,-16'h0099,-16'h0013,16'h0139,16'h00f0,16'h0139,-16'h0058,-16'h0030,16'h00aa,16'h0056,-16'h0057,16'h01a5,16'h001a,16'h0006,16'h00fe,-16'h0085,-16'h0033,16'h0045,-16'h0042,16'h00da,-16'h003f,-16'h0023,-16'h01e0,16'h009e,-16'h007f,-16'h0101,16'h003e,-16'h0087,16'h017b,-16'h00f5,16'h001a,16'h0047,-16'h00a8,-16'h01d0,-16'h0453,16'h00f8,16'h0064,16'h006a,16'h0004,-16'h007d,-16'h00b8,-16'h0004,16'h0174,-16'h000b,-16'h0018,-16'h0086,16'h016a,-16'h00a6,16'h030f,-16'h0077,16'h0289,16'h00e9,16'h00ff,16'h00b4,16'h00c2,16'h0015,-16'h022f,16'h0059,-16'h007c,-16'h0337,-16'h0086,16'h0047,-16'h0041,16'h001c,16'h008b,-16'h0087,-16'h0036,16'h014d,16'h0091,16'h011d,-16'h0048,-16'h007e,16'h0037,16'h0028,-16'h0067,16'h014a,16'h00cd,16'h001c,16'h00fd,-16'h0089,-16'h0038,16'h0027,-16'h0054,16'h014c,16'h0033,-16'h0041,-16'h0204,-16'h001f,-16'h006b,-16'h0180,-16'h0010,-16'h0107,16'h0159,-16'h00dd,16'h000f,16'h00bb,16'h000c,-16'h0217,-16'h03df,16'h0066,-16'h0004,16'h005d,-16'h0089,-16'h0026,-16'h00b2,-16'h0008,16'h0097,-16'h0088,-16'h004e,-16'h0015,16'h0136,-16'h0047,16'h02ce,-16'h0087,16'h0267,16'h00d6,16'h00aa,16'h00fa,16'h00f9,16'h0062,-16'h0330,16'h0097,16'h005d,-16'h029a,-16'h015e,16'h0072,-16'h0058,-16'h0091,16'h00f0,-16'h007c,-16'h00a3,16'h0061,16'h0077,16'h011e,-16'h00cf,-16'h0031,16'h0002,16'h000c,-16'h00cc,16'h0020,16'h0155,16'h003d,16'h000d,-16'h00ad,16'h0035,-16'h005e,-16'h0038,16'h015c,16'h002a,-16'h00f8,-16'h00f0,-16'h0007,-16'h0054,-16'h00e8,16'h007d,-16'h0122,16'h006b,-16'h001c,-16'h0019,16'h011c,16'h0084,-16'h026a,-16'h0230,16'h00bb,16'h0015,16'h0069,-16'h0107,-16'h0041,-16'h00bd,-16'h0030,16'h017c,-16'h00db,-16'h0024,16'h0014,16'h01cf,16'h0047,16'h0308,16'h0015,16'h0259,16'h00af,-16'h0014,16'h0109,16'h0126,16'h0013,-16'h05d7,16'h0003,16'h005e,-16'h02f3,-16'h01e9,16'h0053,-16'h0080,-16'h00cc,16'h00a4,16'h0002,-16'h0104,-16'h004c,16'h00c9,16'h00df,-16'h0038,-16'h0042,16'h000c,-16'h003b,-16'h0055,16'h000c,16'h012e,-16'h00b9,-16'h002b,-16'h0076,16'h0063,-16'h0024,-16'h000b,16'h017b,16'h007c,-16'h00c5,-16'h00ba,-16'h002e,-16'h006a,-16'h005a,-16'h004e,-16'h00d0,16'h0068,-16'h0022,16'h001d,16'h00e6,16'h00d9,-16'h026d,-16'h0095,16'h00a4,-16'h0024,16'h002a,-16'h0066,-16'h0019,-16'h0099,-16'h0050,16'h015f,-16'h00d8,-16'h00c4,16'h0088,16'h0116,16'h0090,16'h02f3,-16'h008e,16'h0296,16'h0127,16'h0058,16'h0111,16'h00ac,-16'h0084,-16'h0516,16'h0080,-16'h0045,-16'h023a,-16'h015e,16'h0043,-16'h0098,-16'h00a9,16'h00d1,16'h0024,-16'h0045,-16'h01c0,16'h00f6,16'h0083,-16'h005c,-16'h0081,-16'h0006,16'h0047,-16'h005e,-16'h0060,16'h00f8,-16'h0084,-16'h0073,-16'h0041,16'h00f9,16'h0000,-16'h0017,16'h01d9,16'h0021,-16'h00ca,-16'h007c,-16'h002c,-16'h0028,16'h0188,-16'h0042,-16'h004f,16'h000b,-16'h005c,-16'h005e,16'h00d4,16'h013b,-16'h0179,16'h0075,16'h0049,-16'h0084,16'h007b,-16'h000b,-16'h0040,-16'h00e1,-16'h0077,16'h0123,-16'h0098,-16'h006f,16'h00c3,-16'h0016,16'h0020,16'h028e,-16'h0129,16'h0257,16'h00ef,16'h0045,16'h00aa,16'h0134,-16'h0033,-16'h03a7,16'h0015,16'h005a,-16'h01fe,-16'h014d,-16'h0053,-16'h005a,-16'h00c7,16'h00e3,16'h0016,-16'h009d,-16'h014c,16'h0104,16'h0049,-16'h003e,-16'h0041,-16'h000b,-16'h0084,16'h0012,-16'h00ce,16'h011f,-16'h0050,-16'h0036,16'h000a,16'h005c,-16'h001f,16'h001a,16'h01cf,-16'h003d,-16'h003e,-16'h005f,-16'h00ac,-16'h0084,16'h018c,-16'h005e,-16'h0080,16'h001c,-16'h0049,-16'h002c,16'h00ab,16'h0163,-16'h0086,16'h00f2,-16'h006c,-16'h0085,16'h007d,-16'h0025,-16'h0016,16'h005f,-16'h0068,16'h012d,-16'h0095,-16'h007d,16'h000c,-16'h00b8,-16'h003a,16'h029d,-16'h0022,16'h0216,16'h013f,16'h009e,16'h0010,16'h0103,16'h000d,-16'h0163,-16'h003b,16'h0077,-16'h022e,-16'h0160,-16'h0016,-16'h003f,-16'h012e,16'h0001,16'h00ad,-16'h00a2,-16'h0123,16'h0141,16'h0043,-16'h003e,-16'h0084,16'h0010,-16'h007e,16'h006e,-16'h007b,16'h00ca,-16'h004b,16'h003c,-16'h000a,16'h002d,-16'h0084,16'h000d,16'h0223,-16'h0023,16'h0028,-16'h00e7,-16'h00c2,16'h001d,16'h01b5,16'h00b7,16'h0036,-16'h000e,-16'h002f,-16'h004c,16'h008f,16'h0161,16'h004d,16'h0128,16'h0069,-16'h006d,16'h00a7,16'h0061,-16'h0018,16'h00e3,-16'h0065,16'h00be,-16'h0147,-16'h00c6,-16'h0079,-16'h00d5,-16'h0064,16'h0262,16'h00a5,16'h020c,16'h01a2,16'h0042,16'h001b,16'h00c3,-16'h002a,-16'h0141,-16'h004e,16'h00e5,-16'h0247,-16'h0166,-16'h0054,16'h0096,-16'h00ed,16'h00da,16'h00ed,-16'h0044,-16'h0063,16'h016d,-16'h00a3,16'h0004,-16'h0040,-16'h0001,-16'h00f3,-16'h0028,-16'h0053,16'h00d4,16'h0060,16'h0056,16'h006f,-16'h0002,-16'h0069,-16'h000e,16'h0215,16'h0043,16'h001b,-16'h007e,-16'h0112,16'h0096,16'h0078,16'h00fb,16'h00bc,16'h0085,-16'h002e,-16'h005f,16'h0075,16'h0162,16'h0155,16'h0122,16'h00ab,-16'h0010,16'h0039,-16'h0012,-16'h000a,16'h0044,-16'h004d,16'h00d4,-16'h0103,-16'h008e,-16'h0046,-16'h00d5,-16'h0075,16'h0202,16'h00dd,16'h0244,16'h027b,16'h006f,-16'h0053,16'h00a5,16'h002e,-16'h0150,-16'h001a,16'h00f6,-16'h01cf,-16'h0158,16'h0063,16'h0044,-16'h012d,16'h00d6,16'h00c7,-16'h0046,16'h00a3,16'h014e,-16'h00c7,-16'h0007,-16'h00f9,-16'h0006,-16'h0092,16'h0001,16'h0014,16'h0117,16'h004c,-16'h0029,-16'h0001,16'h003e,-16'h0032,-16'h0033,16'h016b,16'h0002,16'h0065,16'h00f5,-16'h0081,16'h000e,-16'h01a9,16'h0141,16'h00a4,16'h0034,-16'h000f,-16'h003c,16'h006c,16'h00d4,16'h0102,16'h0156,16'h0096,16'h002f,16'h0058,-16'h000b,-16'h0016,-16'h009e,-16'h0032,16'h00e9,-16'h0045,-16'h007d,-16'h0027,-16'h0040,-16'h00dd,16'h01e2,16'h00d3,16'h0198,16'h0244,16'h0034,-16'h0054,16'h00e5,16'h0073,-16'h01b0,-16'h0033,16'h00e8,-16'h01e1,-16'h0173,16'h0058,-16'h0030,-16'h01c2,16'h0068,16'h0087,16'h002f,16'h0112,16'h0109,-16'h0042,16'h0014,-16'h0071,-16'h001e,-16'h001e,-16'h002d,16'h0008,16'h01b0,16'h00ba,16'h0013,-16'h0016,16'h0064,-16'h0020,-16'h0060,16'h0046,-16'h0012,16'h0103,16'h012c,-16'h00d6,16'h009e,-16'h026c,16'h017e,16'h0174,16'h003c,16'h0017,-16'h0042,16'h0091,-16'h0072,16'h0168,16'h00e0,16'h0091,-16'h0061,16'h0072,16'h0006,16'h0006,-16'h0157,16'h0007,16'h00d1,16'h0076,-16'h00ac,16'h0086,-16'h0023,-16'h0023,16'h01e3,16'h00ef,16'h01b9,16'h023f,-16'h0023,-16'h0094,-16'h0038,16'h011b,-16'h0115,-16'h0124,16'h00db,-16'h01a2,-16'h00d7,16'h00b1,-16'h005b,-16'h01e6,16'h00d1,16'h0102,16'h0010,16'h00e8,16'h0179,-16'h00ab,16'h0082,-16'h008a,-16'h001b,-16'h001c,-16'h0029,-16'h001f,16'h0203,16'h0125,-16'h00cd,-16'h0050,16'h00d8,-16'h005d,16'h0013,-16'h0067,-16'h0078,16'h00bf,16'h0122,-16'h0074,16'h0034,-16'h0167,16'h01b5,16'h01f0,16'h0085,16'h0034,-16'h002c,16'h00ef,-16'h029d,16'h0186,16'h005d,-16'h0057,-16'h0053,-16'h005d,-16'h0022,-16'h0049,-16'h01ac,-16'h001d,-16'h0044,16'h008c,-16'h00b8,16'h0100,16'h0053,16'h00bf,16'h01be,16'h0138,16'h012b,16'h0192,16'h001d,-16'h00ed,-16'h0043,16'h00a1,16'h0003,-16'h0099,16'h00d7,-16'h0173,-16'h0116,16'h00d4,-16'h0093,-16'h0153,16'h0143,16'h018e,-16'h004e,16'h0096,16'h0134,-16'h008b,16'h016d,-16'h00ac,16'h0025,16'h000a,-16'h002e,16'h002d,16'h015e,16'h016e,-16'h00cd,-16'h0039,16'h0051,-16'h016e,16'h0015,-16'h0144,-16'h006e,16'h0077,16'h0145,16'h00ae,-16'h0011,-16'h0091,16'h0156,16'h021b,-16'h000f,16'h0004,-16'h0034,16'h0190,-16'h05f9,16'h015c,16'h000b,-16'h003c,-16'h0022,-16'h0014,-16'h0027,-16'h0099,-16'h00f1,-16'h0025,-16'h0095,16'h009b,16'h002e,16'h0137,-16'h009d,16'h0182,16'h01c9,-16'h006a,16'h017f,16'h014f,-16'h0001,-16'h0095,-16'h0006,-16'h0157,16'h015a,-16'h0112,16'h00ba,-16'h0180,-16'h0142,16'h0112,-16'h003c,-16'h0106,16'h013c,16'h01a1,16'h0021,16'h00d5,16'h0173,-16'h004e,16'h015b,-16'h004e,16'h0031,-16'h001c,16'h0064,16'h0039,16'h01c9,16'h0145,-16'h009c,-16'h0046,16'h00a5,-16'h0148,16'h0019,-16'h01ac,-16'h0009,16'h00a0,16'h0185,16'h011a,16'h0064,-16'h0037,16'h00da,16'h01fb,-16'h00d8,16'h0043,-16'h0033,16'h0179,-16'h07c9,16'h009d,-16'h0038,-16'h0035,-16'h002c,16'h0010,-16'h003d,-16'h00c5,16'h0066,16'h002b,-16'h00fc,16'h0006,16'h00bc,16'h00b4,-16'h00be,16'h0156,16'h0236,-16'h0216,16'h019c,16'h0156,-16'h0034,-16'h0026,-16'h0046,-16'h046c,16'h012e,-16'h00d3,16'h00ce,-16'h0190,-16'h0153,16'h00b3,-16'h0009,-16'h00da,16'h0091,16'h01c2,16'h00db,16'h008a,16'h016c,-16'h0077,16'h0141,16'h001e,16'h001b,16'h0025,16'h007d,-16'h007e,16'h0238,16'h0130,-16'h0126,-16'h0084,16'h00e0,-16'h00b2,-16'h004c,-16'h0294,-16'h0074,16'h0086,16'h01a2,16'h0152,16'h0032,16'h0099,-16'h00a9,16'h01a9,-16'h01f2,16'h0043,-16'h0006,16'h0122,-16'h05ce,-16'h0045,-16'h007b,16'h00d2,-16'h001f,-16'h0033,16'h0043,-16'h010a,16'h01ab,16'h007f,-16'h0167,16'h006e,16'h006b,16'h011c,-16'h00ce,16'h00d7,16'h0140,-16'h0214,16'h00e6,16'h0105,16'h001b,16'h00e7,-16'h0006,-16'h05c1,16'h01b0,-16'h01e7,16'h00d7,-16'h019d,-16'h010a,16'h0043,16'h0043,-16'h00d6,16'h00c9,16'h0171,16'h0103,16'h0095,16'h015b,16'h004b,16'h011c,16'h003b,16'h008e,-16'h008f,16'h00aa,-16'h0002,16'h0266,16'h0100,-16'h0162,-16'h007d,16'h00e8,-16'h00f1,-16'h004b,-16'h02a1,16'h0011,16'h0075,16'h00de,16'h00ac,16'h004f,16'h0014,-16'h02cb,16'h0153,-16'h01b2,-16'h003d,16'h00bd,16'h0076,-16'h02c5,-16'h0077,-16'h0086,16'h00cd,-16'h0064,16'h0022,16'h0169,-16'h00af,16'h01fa,-16'h0037,-16'h0286,16'h001e,16'h0000,16'h0078,-16'h00a5,-16'h005d,16'h0095,-16'h0025,16'h016b,16'h0112,16'h001e,16'h0158,-16'h0082,-16'h056a,16'h0118,-16'h0221,16'h0029,-16'h0174,-16'h002d,16'h009e,-16'h0012,-16'h009b,16'h012d,16'h014f,16'h00ae,-16'h000b,16'h011f,16'h0026,16'h00b8,16'h0031,16'h006b,-16'h003c,16'h0142,-16'h0026,16'h01be,16'h00f1,-16'h00b9,-16'h0051,16'h00a7,-16'h0036,16'h004e,-16'h0329,16'h0054,16'h007b,16'h0060,16'h00c7,16'h011d,-16'h0070,-16'h03f5,16'h015a,-16'h014b,-16'h0022,16'h0034,16'h00d8,-16'h01d3,-16'h003d,-16'h0034,16'h0117,16'h0033,-16'h0008,16'h01d2,-16'h0101,16'h0082,-16'h0033,-16'h02bd,16'h0004,-16'h007a,16'h0095,16'h0027,-16'h012a,16'h011b,16'h0165,16'h0125,16'h0118,16'h0093,16'h0195,-16'h0062,-16'h049a,16'h014c,-16'h0215,-16'h0014,-16'h0174,16'h00db,16'h0089,16'h0000,-16'h00d0,16'h0107,16'h00f8,16'h0053,-16'h006c,16'h0174,-16'h000e,16'h00cb,16'h00ff,16'h0058,16'h0027,16'h0118,16'h0049,16'h0230,16'h0148,-16'h0048,16'h0019,16'h00b8,16'h000e,-16'h0057,-16'h034d,16'h008f,16'h007d,-16'h006c,16'h00f6,16'h00cd,-16'h001d,-16'h02fc,16'h016c,-16'h002f,-16'h0002,16'h0066,16'h00be,-16'h0125,-16'h0053,-16'h00c8,16'h00ab,-16'h0015,-16'h0025,16'h01a3,-16'h011b,-16'h0045,-16'h0073,-16'h02aa,-16'h0071,-16'h0165,16'h0169,16'h003c,-16'h0142,16'h010d,16'h0303,16'h00e3,16'h0117,16'h00b2,16'h0156,-16'h0042,-16'h0378,16'h0104,-16'h0114,-16'h0085,-16'h012d,16'h00e7,16'h0058,-16'h002d,-16'h0026,16'h00ec,16'h00da,16'h00b8,-16'h004c,16'h0208,-16'h004a,16'h0149,16'h013d,16'h0051,-16'h0001,16'h011f,16'h0067,16'h01a3,16'h012f,16'h000d,16'h008f,16'h00d3,16'h0013,16'h0021,-16'h035d,16'h006f,16'h0076,-16'h01a5,16'h0136,16'h00c9,16'h0057,-16'h0139,16'h01d1,16'h0039,16'h001c,16'h0010,16'h00f6,-16'h00cc,16'h0028,-16'h00b2,16'h0007,-16'h00b3,-16'h005c,16'h00cd,-16'h00e4,-16'h00d0,-16'h00d5,-16'h01e6,-16'h000f,-16'h02a5,16'h0082,-16'h009b,-16'h00e1,16'h0182,16'h0387,16'h00ff,16'h0147,16'h00d3,16'h01c0,-16'h000a,-16'h01cb,16'h0109,-16'h006f,-16'h0102,-16'h00ab,16'h00cd,16'h010a,16'h0005,16'h0041,16'h0093,-16'h018a,16'h014e,-16'h0081,16'h026a,16'h0036,16'h01b0,16'h010f,-16'h0082,-16'h004c,16'h00ed,16'h00e9,16'h00b1,16'h0113,16'h0005,16'h00d3,16'h00ef,16'h0116,16'h003d,-16'h0339,-16'h0020,16'h00c1,-16'h0362,16'h015c,16'h0098,-16'h0081,16'h005a,16'h01f7,16'h0170,16'h0046,-16'h0027,16'h006a,-16'h0076,-16'h0051,-16'h00f9,-16'h00b5,-16'h00c1,-16'h004c,16'h00b8,-16'h015d,-16'h01cc,-16'h00cc,-16'h00e2,-16'h0049,-16'h0275,16'h0084,-16'h0087,-16'h000d,16'h01ba,16'h028d,16'h0128,16'h0130,16'h00fd,16'h0164,16'h0009,-16'h011c,16'h00a7,-16'h0055,-16'h00b9,-16'h006d,16'h00b1,16'h016c,-16'h0026,16'h0085,-16'h0058,-16'h027e,16'h0145,-16'h0045,16'h01ce,16'h007c,16'h012b,16'h01c6,-16'h00a0,-16'h00bf,16'h00a8,16'h00a1,16'h003a,16'h007d,-16'h003a,16'h0072,16'h00b9,16'h0114,16'h00d6,-16'h023d,16'h00a2,16'h00fb,-16'h04ab,16'h01de,16'h0077,-16'h0068,16'h0198,16'h01d1,16'h01cc,-16'h0046,-16'h00e8,16'h009a,-16'h0050,-16'h00d4,-16'h0093,-16'h0105,-16'h0048,16'h004d,16'h008b,-16'h00ac,-16'h021f,16'h00fb,-16'h0086,16'h0052,-16'h02cd,16'h008b,-16'h006b,-16'h004c,16'h02d5,16'h012b,16'h0054,16'h00a7,16'h00fd,16'h01c4,16'h003b,-16'h0132,16'h014c,16'h0053,16'h000c,-16'h0087,16'h00b8,16'h0193,-16'h0075,-16'h0083,-16'h0146,-16'h031a,16'h013e,-16'h0033,16'h00fb,16'h0043,-16'h00a1,16'h01dc,-16'h0068,-16'h0078,-16'h0025,16'h007d,-16'h001a,16'h0113,-16'h0036,16'h00ca,16'h00b5,16'h0148,16'h0055,-16'h0202,16'h008a,16'h00a5,-16'h0414,16'h00ca,16'h0050,16'h0041,16'h01d2,16'h01ae,16'h01ba,16'h007c,-16'h00e1,16'h0085,-16'h0026,-16'h0114,-16'h0115,-16'h00ba,-16'h003e,16'h0084,16'h009c,-16'h005d,-16'h013a,16'h00b2,-16'h009f,-16'h0012,-16'h01f6,16'h00a2,-16'h004f,-16'h0059,16'h02c3,16'h007b,16'h0041,16'h007a,16'h01cf,16'h01cb,16'h00e2,-16'h00e9,16'h0124,16'h011b,-16'h004c,-16'h003e,16'h013e,16'h01e7,-16'h00d6,-16'h001d,-16'h00bd,-16'h0209,16'h010b,16'h003f,16'h00dc,16'h001c,-16'h01a4,16'h01e6,16'h0037,-16'h0038,-16'h0022,-16'h000f,-16'h0104,-16'h020d,-16'h0001,-16'h001b,16'h0010,16'h0071,16'h028e,-16'h014f,16'h00d6,16'h003e,16'h0069,16'h00c7,16'h0014,-16'h01f8,16'h00dc,16'h01bf,-16'h0017,-16'h005b,-16'h0016,16'h0121,-16'h0119,16'h0000,16'h02dc,16'h0154,-16'h00a4,16'h0121,16'h00ab,-16'h00b5,16'h00b6,16'h00b5,-16'h00d7,-16'h005b,16'h004b,-16'h000a,-16'h0098,16'h007c,16'h0083,16'h01a7,16'h0136,16'h00ae,-16'h00b8,16'h0154,16'h0041,16'h01ad,-16'h0127,-16'h00c5,16'h0116,-16'h001d,16'h0065,-16'h01eb,-16'h00b8,-16'h010b,-16'h0068,-16'h0019,16'h0144,-16'h0098,16'h00de,16'h000b,16'h0099,-16'h00b7,16'h008a,-16'h00d8,-16'h0021,16'h00b3,-16'h0148,-16'h0116,-16'h0001,-16'h0096,16'h006d,16'h0037,16'h0210,-16'h0224,16'h014c,16'h00c6,-16'h0059,16'h006a,16'h0061,-16'h0105,16'h00a2,16'h011b,16'h0004,-16'h0036,-16'h00b9,16'h00c0,-16'h00d5,-16'h006c,16'h029c,16'h00e2,16'h002b,16'h01c4,16'h0003,-16'h0072,16'h0036,16'h0010,-16'h00ee,-16'h007b,16'h007b,-16'h004c,-16'h00d1,16'h0040,16'h0051,16'h00bf,16'h017d,16'h00ad,-16'h015c,16'h0101,16'h0015,16'h0165,-16'h0122,-16'h003d,16'h0146,-16'h00b4,16'h0152,-16'h022f,-16'h016b,-16'h00b4,-16'h0019,16'h0038,16'h0110,16'h0032,16'h00cd,16'h0029,16'h0032,-16'h0054,16'h0069,-16'h0090,-16'h009b,16'h0105,-16'h01f6,-16'h00a7,16'h001f,-16'h00fe,16'h0030,16'h0049,16'h011d,-16'h0230,16'h00ac,16'h01a0,-16'h0174,16'h014b,-16'h002a,16'h006c,16'h006b,16'h0088,-16'h0011,-16'h0074,-16'h006a,16'h007d,-16'h0102,-16'h0032,16'h01b2,16'h00c3,-16'h0073,16'h0228,16'h0020,-16'h00fc,-16'h00a2,16'h008a,-16'h0077,-16'h006c,16'h0060,-16'h0047,-16'h00df,-16'h00b8,16'h0026,16'h00a0,16'h0256,16'h005b,-16'h019a,16'h00ab,16'h0024,16'h0119,-16'h01e4,16'h0039,16'h00da,-16'h0065,16'h01f6,-16'h0180,-16'h00d7,-16'h00ad,16'h00b0,-16'h0069,16'h00dd,16'h0063,16'h0106,16'h0027,-16'h006b,-16'h0084,16'h0096,-16'h00a8,-16'h010e,16'h01a2,-16'h0291,-16'h0008,16'h004f,-16'h00a4,-16'h0033,16'h00db,16'h008e,-16'h017b,16'h0031,16'h012b,-16'h016d,16'h00cb,16'h004d,16'h00fd,16'h0005,16'h005e,16'h0039,-16'h0028,-16'h00da,16'h0124,-16'h005a,-16'h0049,16'h00ba,16'h004f,-16'h0010,16'h0225,-16'h004a,-16'h0028,-16'h00b7,-16'h000c,16'h006e,-16'h004b,16'h0037,-16'h008a,-16'h00bc,-16'h0064,16'h012e,16'h001f,16'h021a,16'h00bd,-16'h0169,16'h00ab,16'h005d,16'h00fb,-16'h01e6,16'h0010,16'h00a2,-16'h00d3,16'h0255,-16'h0106,-16'h0113,16'h0024,-16'h000f,16'h0000,16'h012f,16'h00bc,16'h0068,16'h00fc,16'h002a,-16'h0047,16'h0116,-16'h010d,-16'h0125,16'h01d7,-16'h031a,16'h009e,-16'h000d,-16'h0048,16'h0009,16'h0097,16'h0024,-16'h00eb,-16'h008c,16'h00c4,-16'h01e8,16'h0159,-16'h0066,16'h00d9,-16'h00b1,16'h001b,16'h007e,-16'h001c,-16'h00bc,16'h00f1,-16'h0013,-16'h008f,-16'h00e2,16'h0044,-16'h0097,16'h0105,-16'h00a6,16'h0037,-16'h0082,16'h0008,16'h0107,-16'h0043,-16'h003f,-16'h00b9,-16'h00f3,16'h0047,16'h01ca,16'h000f,16'h0279,16'h010b,-16'h006a,16'h011b,16'h00ba,16'h00db,-16'h01d8,16'h0069,16'h00c0,-16'h014e,16'h025b,-16'h0033,-16'h009b,16'h00f1,16'h0061,16'h0007,16'h0097,16'h0152,16'h00b4,16'h00e7,-16'h0036,-16'h0045,16'h0166,-16'h0099,-16'h00f1,16'h01b5,-16'h01c2,16'h008d,-16'h00ad,-16'h00e4,16'h002e,16'h00c8,-16'h0003,-16'h005c,16'h0011,16'h005f,-16'h0158,16'h00cf,-16'h0035,16'h0039,-16'h0072,16'h0018,16'h0019,-16'h0080,-16'h0047,16'h00cc,-16'h0055,-16'h00fc,-16'h0293,16'h00c4,16'h0035,16'h0181,-16'h0031,16'h0049,-16'h0005,-16'h002a,16'h0179,16'h0055,16'h00ba,-16'h0100,16'h0041,16'h0020,16'h0217,16'h0030,16'h0298,16'h00d2,16'h005d,16'h008b,16'h0033,16'h00d1,-16'h022c,16'h00b7,16'h001e,-16'h01a4,16'h01ac,-16'h0061,-16'h006e,16'h0129,16'h0089,-16'h009c,16'h0052,16'h00c1,16'h00c8,16'h00d4,-16'h001b,-16'h0026,16'h012a,-16'h00d6,-16'h00a5,16'h01f3,-16'h0065,16'h0023,-16'h0115,-16'h00e8,16'h004c,16'h00d5,-16'h0018,16'h00ca,-16'h0035,16'h0016,-16'h0175,16'h00a4,-16'h0092,-16'h00bb,-16'h006d,-16'h0064,16'h002e,-16'h0146,-16'h0089,16'h0098,-16'h0100,-16'h0147,-16'h0426,16'h0112,-16'h003e,16'h00f6,16'h0008,-16'h0022,-16'h0046,-16'h002b,16'h011c,-16'h0027,16'h0099,-16'h00b8,16'h0120,-16'h0026,16'h0241,16'h0000,16'h02ea,16'h0092,16'h00a1,16'h00c9,16'h00a0,16'h0118,-16'h0267,16'h0092,-16'h002a,-16'h0232,16'h00df,-16'h002a,-16'h004d,16'h00c7,16'h0059,-16'h00a7,-16'h002c,16'h017c,16'h00c4,16'h015f,-16'h006d,-16'h009b,16'h0142,-16'h0026,-16'h00c3,16'h010e,16'h009e,16'h002d,-16'h00f4,-16'h00aa,16'h001d,16'h0061,16'h001e,16'h01df,-16'h0059,16'h003c,-16'h01da,16'h009b,-16'h00f9,-16'h01e0,-16'h0048,-16'h004b,16'h0080,-16'h00ba,-16'h0016,16'h0119,-16'h00d5,-16'h011d,-16'h04d3,16'h00f7,-16'h0079,16'h0148,-16'h0026,-16'h0022,-16'h0053,-16'h0095,16'h012c,16'h0029,-16'h002b,-16'h0065,16'h0092,-16'h004c,16'h0299,-16'h0002,16'h029e,16'h001d,16'h00b6,16'h010f,16'h0088,16'h00e5,-16'h0363,16'h0021,16'h0051,-16'h020e,-16'h00bc,-16'h0049,-16'h00f6,16'h012c,16'h0093,-16'h002d,-16'h00c7,16'h0083,16'h00b5,16'h00ef,-16'h0052,-16'h009c,16'h00ff,-16'h0047,-16'h00d4,16'h008d,16'h01a8,-16'h003b,-16'h0230,-16'h0086,-16'h005e,-16'h004f,-16'h002a,16'h01f5,-16'h009c,16'h0037,-16'h0199,16'h006c,-16'h00a0,-16'h01f8,16'h000a,-16'h0045,16'h00f0,-16'h007f,16'h001e,16'h0066,-16'h006d,-16'h0266,-16'h02a4,16'h0115,16'h000e,16'h00ed,-16'h0054,-16'h0005,-16'h00ab,-16'h0061,16'h014b,-16'h00c6,16'h000b,-16'h0031,16'h00c7,16'h005c,16'h029c,-16'h009a,16'h029d,16'h0000,16'h00a0,16'h00c7,16'h000e,16'h0069,-16'h0538,-16'h002e,16'h0024,-16'h009e,-16'h0148,16'h0019,-16'h0045,16'h00a8,16'h00c9,16'h003c,-16'h0125,-16'h00eb,16'h00a0,16'h00ad,-16'h00d1,-16'h0095,16'h00d0,-16'h0015,-16'h0072,16'h00ff,16'h011b,-16'h003a,-16'h024c,-16'h002a,-16'h0093,-16'h0015,-16'h0017,16'h0293,-16'h0063,-16'h0038,-16'h00b4,16'h0099,-16'h0059,-16'h00dc,-16'h0031,-16'h007a,16'h009e,-16'h001b,16'h0010,16'h0133,16'h0076,-16'h02d4,-16'h00a4,16'h00ee,-16'h000d,16'h007f,16'h0007,-16'h0070,-16'h0177,-16'h000e,16'h01a1,-16'h0071,-16'h00a2,16'h0024,16'h014c,16'h0097,16'h035a,-16'h003b,16'h02c1,16'h002e,-16'h0023,16'h0146,16'h009d,-16'h0011,-16'h055f,16'h000c,16'h008f,-16'h0066,-16'h01b5,-16'h0071,-16'h0025,16'h0065,16'h00b4,16'h000d,-16'h0190,-16'h01c9,16'h00b1,16'h00b8,-16'h00b4,-16'h0037,16'h0048,16'h000c,-16'h00ad,16'h0030,16'h0089,-16'h00d1,-16'h01b7,-16'h0061,-16'h004b,-16'h0003,-16'h0050,16'h029d,-16'h0024,16'h0000,-16'h00d8,16'h0050,-16'h00c0,16'h00e1,-16'h00aa,16'h0002,-16'h0025,-16'h0043,16'h0025,16'h0105,16'h00bc,-16'h02be,16'h0049,16'h00a0,16'h0023,16'h00fb,-16'h0011,-16'h0062,-16'h0135,-16'h002e,16'h01a3,16'h0011,-16'h0102,16'h00a9,16'h007a,16'h0006,16'h033b,-16'h0088,16'h0241,16'h0116,16'h003b,16'h010d,16'h00e8,16'h0088,-16'h0413,-16'h0020,16'h0014,-16'h00d8,-16'h01d0,-16'h0036,16'h000c,16'h00b2,16'h0112,16'h002d,-16'h0120,-16'h01d9,16'h00cb,16'h001f,-16'h00a1,-16'h00b2,16'h00c9,-16'h0032,-16'h007c,-16'h008c,16'h009f,-16'h007e,-16'h020f,16'h0007,-16'h0077,16'h0014,16'h0034,16'h01ee,16'h0040,-16'h00a0,-16'h0068,16'h00d2,-16'h0093,16'h020d,-16'h0132,16'h0019,-16'h0070,16'h0016,-16'h0007,16'h00f9,16'h013d,-16'h0146,16'h008b,-16'h0024,-16'h00eb,16'h00c5,16'h0060,-16'h0008,-16'h0071,16'h0057,16'h016e,-16'h0041,-16'h00f6,16'h004a,-16'h00cd,16'h0039,16'h0369,-16'h010e,16'h0258,16'h00ce,16'h008d,16'h00ee,16'h00bd,16'h0098,-16'h0298,-16'h001b,16'h008d,-16'h00c1,-16'h01de,-16'h003a,-16'h0060,16'h0042,16'h010b,-16'h0070,-16'h013b,-16'h0165,16'h015e,16'h004a,-16'h0026,-16'h008d,16'h0029,-16'h0077,16'h001c,-16'h006f,16'h00c1,-16'h0024,-16'h0289,16'h0013,-16'h0014,-16'h002e,16'h00c1,16'h0211,16'h002e,-16'h0040,-16'h00a5,16'h002c,-16'h0044,16'h01f4,-16'h00e0,-16'h0012,-16'h001e,-16'h001a,16'h003f,16'h00ee,16'h01e4,-16'h0007,16'h013d,-16'h0043,-16'h0042,16'h013f,-16'h002f,-16'h0006,-16'h0023,16'h001b,16'h01ac,-16'h00b3,-16'h00bc,16'h003a,-16'h0202,16'h005b,16'h0313,-16'h0002,16'h023b,16'h00ae,16'h002c,16'h0054,16'h0092,16'h0023,-16'h0099,-16'h0083,16'h0124,-16'h00c0,-16'h0221,-16'h0086,16'h004f,16'h008a,16'h00c0,16'h0048,-16'h0103,-16'h0018,16'h01e4,-16'h003f,16'h0025,-16'h003c,-16'h0065,-16'h001a,-16'h0057,-16'h005d,16'h00b2,16'h005a,-16'h0219,16'h004a,16'h001f,-16'h0003,16'h002f,16'h01c0,-16'h0008,16'h0018,-16'h00e0,-16'h00b6,-16'h00ad,16'h0120,16'h0047,16'h00c2,-16'h0067,-16'h0038,16'h000a,16'h007c,16'h020e,16'h0170,16'h00a3,16'h005c,-16'h0020,16'h00d2,16'h003e,-16'h0090,16'h009e,-16'h003b,16'h013d,-16'h00cf,-16'h0116,-16'h006d,-16'h01b8,-16'h0002,16'h02db,16'h005a,16'h0255,16'h00dc,16'h0034,16'h009b,16'h00ca,16'h00b9,-16'h010e,-16'h0013,16'h007d,-16'h0134,-16'h0237,-16'h000a,16'h0052,-16'h0008,16'h0122,16'h0088,-16'h00cd,16'h008f,16'h01d8,-16'h00ae,16'h0063,16'h0030,16'h000a,-16'h00aa,-16'h0037,-16'h003e,16'h010f,16'h00d2,-16'h021e,-16'h0023,-16'h005d,16'h0042,16'h002f,16'h0113,16'h0019,16'h0038,-16'h00a9,-16'h00d3,16'h000b,-16'h00d7,16'h0119,16'h015f,16'h005c,16'h0025,-16'h0028,16'h003c,16'h029d,16'h018b,16'h013e,16'h0076,16'h001c,16'h00c2,16'h0029,16'h0046,16'h002a,-16'h0074,16'h016d,-16'h004e,-16'h0123,-16'h00e4,-16'h007a,-16'h008d,16'h020f,16'h00a9,16'h0259,16'h0155,-16'h001a,16'h0052,16'h00fd,16'h004e,-16'h0166,-16'h0060,16'h00e2,-16'h0013,-16'h0184,16'h007f,16'h005e,-16'h0062,16'h00fa,16'h0045,-16'h005e,16'h014f,16'h01a1,-16'h00a7,16'h0064,-16'h0018,16'h007b,-16'h0075,16'h003e,-16'h001e,16'h01b2,16'h0171,-16'h01e9,16'h0056,16'h0062,16'h0011,-16'h000a,-16'h0010,-16'h006a,16'h0052,16'h00bd,-16'h00ca,16'h004f,-16'h01a0,16'h0133,16'h011f,16'h006f,-16'h000f,16'h0015,16'h003b,16'h01a7,16'h017b,16'h00dc,16'h005c,-16'h002c,16'h0105,16'h0042,-16'h0030,-16'h008c,-16'h001f,16'h00bb,16'h0083,-16'h0083,16'h0007,-16'h000e,-16'h011f,16'h01d0,16'h0121,16'h0247,16'h018a,16'h0042,16'h0036,16'h0073,16'h010e,-16'h00f5,16'h000f,16'h00ca,-16'h001b,-16'h004a,16'h0104,16'h0092,-16'h0064,16'h0103,16'h00ef,-16'h00e3,16'h016c,16'h01aa,-16'h00f3,16'h0046,-16'h003c,-16'h001c,-16'h004d,-16'h000c,16'h004b,16'h01df,16'h0186,-16'h02b1,16'h0060,16'h00ad,-16'h0038,16'h0059,-16'h0054,16'h0023,16'h0090,16'h0184,-16'h008d,16'h0095,-16'h026c,16'h0204,16'h018e,-16'h0019,16'h008d,-16'h0009,16'h0097,16'h0056,16'h010c,16'h009b,16'h00ba,-16'h00a1,16'h0100,16'h0076,-16'h003c,-16'h024d,16'h0043,16'h0029,16'h00a9,-16'h009a,16'h005e,16'h005f,-16'h00e0,16'h01a0,16'h00e8,16'h01c5,16'h0174,16'h0008,-16'h0082,16'h008a,16'h018d,-16'h00d5,-16'h00ba,16'h00b4,16'h009a,-16'h014e,16'h0135,16'h007a,-16'h006d,16'h0114,16'h014a,-16'h0123,16'h0052,16'h016b,-16'h0090,16'h001a,-16'h0019,-16'h002c,-16'h003a,-16'h00af,16'h0024,16'h01bd,16'h017e,-16'h02a9,16'h003d,16'h005d,16'h0013,16'h001c,-16'h0171,-16'h0099,16'h00b6,16'h01a3,-16'h0070,16'h0113,-16'h00b3,16'h0239,16'h0255,-16'h003a,16'h00b3,-16'h00af,16'h00f5,-16'h0224,16'h018e,16'h0066,16'h0019,-16'h0036,16'h0096,16'h0049,-16'h0086,-16'h022c,-16'h0011,-16'h00a9,16'h004f,-16'h0055,16'h00d3,-16'h0034,16'h0050,16'h01b1,16'h00de,16'h0199,16'h0101,-16'h001d,-16'h006c,16'h0023,16'h0129,16'h0081,-16'h0093,16'h00dc,16'h0083,-16'h0124,16'h0178,16'h000b,-16'h00e8,16'h00d4,16'h0126,-16'h00ef,16'h0031,16'h0146,16'h0003,16'h011f,-16'h00c7,16'h0014,-16'h004b,-16'h009f,16'h003b,16'h017f,16'h0167,-16'h0296,-16'h002a,16'h00ea,-16'h00b8,16'h0017,-16'h01ff,-16'h0041,16'h0052,16'h011b,16'h001d,16'h0094,-16'h00a8,16'h01d6,16'h0261,-16'h0037,16'h001f,-16'h0022,16'h016a,-16'h0664,16'h00a1,-16'h001a,-16'h0012,-16'h0019,16'h0050,16'h002f,-16'h007f,-16'h0184,16'h0021,-16'h00fe,16'h0081,16'h0012,16'h00c9,-16'h00ec,16'h0111,16'h0155,16'h000d,16'h0183,16'h008d,-16'h0031,-16'h0045,16'h00ac,16'h0052,16'h00e4,-16'h0064,16'h00af,16'h000b,-16'h01a2,16'h018f,-16'h0013,-16'h009b,16'h0104,16'h0111,-16'h003d,16'h002d,16'h0160,16'h003d,16'h0167,-16'h0055,16'h002d,-16'h0059,16'h006a,16'h001b,16'h01a8,16'h0172,-16'h024e,-16'h0073,16'h00e6,-16'h0082,16'h0065,-16'h024a,-16'h0037,-16'h00ab,16'h01a5,16'h00b2,16'h004f,16'h0032,16'h00cf,16'h0257,-16'h00d7,16'h003b,-16'h0064,16'h0159,-16'h090d,16'h0026,16'h0021,16'h0042,-16'h0035,16'h0040,16'h004d,-16'h00a9,16'h0032,16'h007a,-16'h0121,16'h0081,16'h005f,16'h016a,-16'h0119,16'h0201,16'h0180,-16'h0271,16'h0190,-16'h0068,16'h0020,-16'h0016,16'h0050,-16'h022b,16'h013a,16'h0011,16'h00b9,16'h0062,-16'h0135,16'h00b3,-16'h001c,-16'h00bb,16'h00eb,16'h00dc,16'h0085,16'h0049,16'h0162,-16'h007c,16'h0163,-16'h0038,16'h0017,-16'h0074,16'h0083,-16'h009b,16'h0177,16'h0174,-16'h0287,-16'h0094,16'h00e8,-16'h00af,-16'h0001,-16'h0284,16'h000a,-16'h001e,16'h01bb,16'h00e5,16'h0011,16'h003a,-16'h010b,16'h018d,-16'h0169,-16'h0013,-16'h0063,16'h015a,-16'h065a,16'h0003,-16'h000c,16'h00da,-16'h0071,16'h0039,16'h00b5,-16'h0144,16'h01d0,16'h0007,-16'h0176,16'h0083,16'h00ba,16'h0108,-16'h0094,16'h00e3,16'h01a8,-16'h02b0,16'h01d7,-16'h0001,-16'h005b,16'h010d,16'h004c,-16'h05c9,16'h00fe,-16'h0048,16'h00bb,-16'h0002,-16'h0089,16'h0066,16'h000b,-16'h00f2,16'h011f,16'h0112,16'h0110,-16'h003f,16'h019d,16'h000b,16'h00ed,-16'h0030,16'h00b2,16'h0037,16'h00e7,16'h004b,16'h012d,16'h019a,-16'h02cf,-16'h0087,16'h00d0,-16'h006f,16'h0001,-16'h02b7,-16'h0013,-16'h0044,16'h00c5,16'h00be,16'h0069,-16'h003a,-16'h02b5,16'h0152,-16'h0294,16'h0027,-16'h0026,16'h00d4,-16'h02a1,-16'h0050,16'h0087,16'h0158,-16'h0026,-16'h0057,16'h0190,-16'h0070,16'h0210,16'h001c,-16'h02a3,16'h0008,16'h00dd,16'h008c,16'h0021,-16'h00c8,16'h011c,-16'h0112,16'h0154,16'h0044,16'h009f,16'h017e,-16'h0001,-16'h06d4,16'h018c,-16'h011c,-16'h0067,-16'h000d,16'h0068,16'h0056,16'h000c,16'h0000,16'h01bc,16'h00b0,16'h00fc,-16'h0098,16'h017f,16'h004e,16'h0109,16'h0016,16'h00ab,16'h0042,16'h0169,16'h002b,16'h00f0,16'h01a8,-16'h0314,-16'h008e,16'h002c,16'h001f,-16'h001b,-16'h027b,16'h0048,16'h0047,16'h00b3,16'h0056,16'h0086,-16'h003d,-16'h04d0,16'h019c,-16'h0195,16'h000f,16'h001e,16'h00f0,-16'h0171,-16'h00a1,-16'h0044,16'h00d9,16'h0007,16'h0012,16'h01d4,-16'h00b8,16'h00c1,-16'h0036,-16'h02db,-16'h0071,-16'h0048,16'h00bf,16'h003b,-16'h0163,16'h00b1,16'h017b,16'h0160,-16'h001e,16'h006e,16'h0191,16'h0007,-16'h0629,16'h0163,-16'h00fd,-16'h004f,16'h0038,16'h007c,16'h00c5,-16'h004c,-16'h00a9,16'h0184,16'h00db,16'h00e8,-16'h0085,16'h0200,-16'h001c,16'h00b5,16'h0098,16'h00b2,16'h0053,16'h0135,16'h0056,16'h00c3,16'h01f9,-16'h0290,-16'h0072,16'h00dc,16'h007e,16'h009c,-16'h02d9,16'h0001,16'h0075,-16'h00a8,16'h0085,16'h00ea,-16'h0095,-16'h03ec,16'h01da,-16'h001c,-16'h001b,16'h0051,16'h00a9,-16'h0125,16'h0008,16'h0005,16'h008b,-16'h0020,-16'h0068,16'h024c,-16'h00ed,-16'h0035,-16'h006d,-16'h027d,-16'h007b,-16'h0126,16'h011d,16'h0071,-16'h0177,16'h0167,16'h02e2,16'h0123,16'h002c,16'h0083,16'h0180,-16'h002f,-16'h04da,16'h0101,-16'h0033,-16'h006c,-16'h0008,16'h00e9,16'h00b6,-16'h012c,-16'h003b,16'h0122,-16'h0031,16'h0111,-16'h00e5,16'h025d,-16'h0004,16'h0157,16'h00fc,16'h0057,16'h003a,16'h00e0,16'h005f,16'h00b7,16'h016e,-16'h0133,-16'h001e,16'h0086,16'h0075,16'h0028,-16'h0322,16'h0038,16'h00b0,-16'h00f0,16'h00e7,16'h004e,-16'h009b,-16'h0214,16'h017b,16'h00ac,16'h0066,16'h000e,16'h00af,-16'h00a2,16'h0046,16'h0050,16'h00b7,-16'h00b1,-16'h00ef,16'h014d,-16'h00ef,-16'h0107,-16'h0133,-16'h0196,-16'h00a0,-16'h0287,16'h00cc,-16'h0034,-16'h0105,16'h018f,16'h035f,16'h00ed,16'h0063,16'h00b2,16'h019e,16'h0045,-16'h0321,16'h00a5,16'h0035,-16'h006f,16'h0005,16'h00d4,16'h0178,-16'h0110,16'h002a,16'h0114,-16'h01c6,16'h0137,-16'h0063,16'h01f6,-16'h0025,16'h0197,16'h0139,-16'h0062,-16'h003e,16'h000b,16'h009f,16'h0000,16'h011b,-16'h00dc,16'h0010,16'h0070,16'h0118,16'h0081,-16'h02d3,16'h0018,16'h0078,-16'h02b7,16'h0137,16'h0007,-16'h005e,16'h0048,16'h014a,16'h0121,16'h00d4,-16'h0043,16'h0072,-16'h0089,-16'h0052,-16'h007f,16'h0009,-16'h00a9,16'h0006,16'h00d2,-16'h0098,-16'h0185,-16'h00e0,-16'h013e,-16'h00c4,-16'h0241,16'h00b9,-16'h0127,16'h003b,16'h0245,16'h02af,16'h00dc,16'h008b,16'h00f4,16'h0215,-16'h001a,-16'h01d3,16'h00a2,-16'h007f,16'h0051,16'h0044,16'h00a4,16'h014a,-16'h0064,-16'h0001,-16'h0030,-16'h0321,16'h01d3,-16'h009c,16'h016c,16'h0051,16'h0039,16'h018b,-16'h002d,-16'h00a8,16'h000d,16'h002e,-16'h00ab,16'h00a4,-16'h00d3,16'h0080,-16'h0021,16'h0145,16'h0124,-16'h0255,16'h003b,16'h0102,-16'h03f5,16'h0156,16'h0076,-16'h0055,16'h0227,16'h010e,16'h01ab,16'h005d,-16'h0018,16'h00a1,-16'h00a9,-16'h00fc,-16'h0025,-16'h009c,-16'h0102,16'h0031,16'h00bf,-16'h00c2,-16'h01e6,16'h0047,-16'h0095,16'h004c,-16'h0258,16'h00a8,-16'h010b,16'h003c,16'h0297,16'h012b,16'h0081,16'h006a,16'h0149,16'h0232,16'h00bc,-16'h0167,16'h009f,-16'h003c,16'h0014,16'h0006,16'h0073,16'h01cf,-16'h0047,-16'h0026,-16'h00d6,-16'h02f6,16'h01df,-16'h0071,16'h0151,-16'h001f,-16'h010d,16'h01ac,-16'h0092,-16'h0058,16'h0028,16'h0077,-16'h0086,16'h000a,-16'h0060,16'h0029,-16'h005d,16'h0194,16'h00e1,-16'h01ba,16'h0027,16'h0070,-16'h04d1,16'h0120,16'h001c,-16'h004c,16'h0217,16'h0162,16'h01f1,16'h005b,-16'h0045,16'h00e9,-16'h0005,-16'h00bf,-16'h00ba,-16'h007a,-16'h00ba,16'h00e5,16'h0095,-16'h0068,-16'h0180,16'h00d6,-16'h007e,16'h0026,-16'h0244,16'h0095,-16'h007d,16'h0000,16'h033f,16'h0072,16'h00ee,16'h007b,16'h017b,16'h022b,16'h00dc,-16'h010a,16'h00fc,16'h0088,16'h005d,16'h0027,16'h00f7,16'h01b7,-16'h00c9,-16'h0042,-16'h00d5,-16'h025e,16'h0108,16'h003e,16'h0125,-16'h002e,-16'h01fc,16'h020f,16'h0085,-16'h0086,16'h0038,16'h00f6,-16'h0152,-16'h0188,-16'h0097,-16'h0064,-16'h0034,16'h0097,16'h026b,-16'h01ac,16'h0168,16'h00c0,16'h0036,16'h00c1,16'h0062,-16'h00ad,16'h00f1,16'h013f,-16'h016f,-16'h00a7,-16'h0050,16'h00d0,-16'h0155,16'h002a,16'h0209,16'h00ec,-16'h000d,16'h01a4,16'h00a8,-16'h009e,16'h006e,16'h00d2,-16'h00cf,-16'h0053,16'h0098,-16'h0033,-16'h0008,16'h003a,16'h0029,16'h01ac,16'h012f,16'h00b7,-16'h0135,16'h00ff,-16'h0008,16'h011d,-16'h00e4,-16'h00d1,16'h015a,-16'h0067,16'h0034,-16'h017c,-16'h004c,-16'h0107,-16'h0020,16'h000f,16'h00d7,16'h0007,16'h01be,16'h005a,16'h001a,-16'h00a8,16'h00a1,16'h0009,16'h0018,16'h00cb,-16'h0189,-16'h00d6,-16'h0054,-16'h000f,16'h004a,16'h0046,16'h01c6,-16'h0202,16'h00a3,16'h00f4,-16'h0043,16'h00bf,-16'h000e,-16'h0057,16'h00d5,16'h00fd,-16'h010e,-16'h006d,-16'h006a,16'h0086,-16'h007f,-16'h0011,16'h0228,16'h00c4,16'h000d,16'h01ee,16'h00b7,-16'h00df,16'h0005,16'h00d2,-16'h00f2,16'h0021,16'h006e,-16'h0041,-16'h008f,-16'h005e,-16'h001c,16'h00da,16'h01b9,16'h00b2,-16'h0182,16'h00dd,-16'h0070,16'h0173,-16'h0192,-16'h0065,16'h0091,-16'h0055,16'h019b,-16'h007a,-16'h0134,-16'h00d2,16'h0054,-16'h0028,16'h010a,16'h00b3,16'h011e,16'h00aa,16'h002d,16'h0002,16'h0088,-16'h0029,-16'h006a,16'h00d2,-16'h0250,-16'h0040,-16'h00cc,16'h0043,16'h0074,16'h007c,16'h00ed,-16'h0250,16'h0020,16'h01d1,-16'h0147,16'h0156,-16'h0031,16'h00c7,-16'h002d,16'h00b3,-16'h0039,-16'h0031,-16'h00db,16'h007b,-16'h0021,-16'h00c7,16'h013b,16'h005e,-16'h002c,16'h021a,16'h0016,-16'h0064,-16'h00ef,16'h00aa,-16'h0078,-16'h0034,-16'h0027,-16'h0080,-16'h010d,-16'h00bb,16'h0016,16'h003d,16'h01d2,16'h00c5,-16'h015d,16'h0012,16'h0062,16'h013b,-16'h0235,-16'h004c,16'h00c9,-16'h0056,16'h01d3,16'h0033,-16'h0107,-16'h005e,16'h002f,-16'h000b,16'h00da,16'h015a,16'h0085,16'h0062,16'h004f,-16'h002c,16'h00cc,-16'h0031,-16'h0122,16'h0113,-16'h0307,16'h0010,-16'h00ef,-16'h0046,16'h000b,16'h00f2,-16'h0018,-16'h01c7,-16'h006b,16'h0141,-16'h00db,16'h00ed,-16'h005c,16'h0154,-16'h0087,16'h0004,-16'h00b0,-16'h0084,-16'h00e5,16'h001b,-16'h0092,-16'h00f3,16'h00b8,16'h006a,-16'h0071,16'h024a,16'h0040,-16'h0073,-16'h0083,16'h009e,-16'h000b,16'h0029,16'h0000,-16'h0111,-16'h00f3,-16'h004d,16'h0015,-16'h008e,16'h0214,16'h010c,-16'h0134,16'h002f,-16'h0022,16'h013d,-16'h022f,-16'h0065,16'h00ff,-16'h0069,16'h020b,-16'h000a,-16'h010b,-16'h003d,16'h007a,-16'h0021,16'h0091,16'h0104,16'h003d,16'h00c7,-16'h004d,16'h0002,16'h013d,-16'h00c7,-16'h010a,16'h0177,-16'h022e,16'h007a,-16'h01d2,16'h001d,16'h0044,16'h00e0,16'h0088,-16'h013b,-16'h004c,16'h015e,-16'h00b1,16'h0150,-16'h0039,16'h00b0,-16'h00fa,16'h0075,-16'h00eb,-16'h0030,-16'h0133,16'h00f3,-16'h0077,-16'h0056,-16'h0142,16'h00a4,-16'h0014,16'h015d,16'h0080,16'h003e,16'h005a,16'h001e,16'h00a0,-16'h0012,16'h0027,-16'h00b3,-16'h0076,16'h0029,16'h0093,-16'h004e,16'h023e,16'h011a,-16'h0078,16'h00bb,16'h0092,16'h014e,-16'h02ae,16'h000b,16'h00e7,-16'h0025,16'h0287,16'h0032,-16'h00ec,16'h0089,16'h00de,-16'h0005,16'h009b,16'h0141,16'h003f,16'h00f6,-16'h0008,-16'h0071,16'h017f,-16'h00c1,-16'h0074,16'h0100,-16'h0131,-16'h0002,-16'h01ee,16'h0007,16'h006e,16'h0150,16'h0036,-16'h0024,-16'h00b3,16'h006c,-16'h008a,16'h012b,-16'h00d2,-16'h000a,-16'h0079,16'h0080,-16'h0198,-16'h0076,-16'h0130,16'h005f,-16'h009f,-16'h0089,-16'h02ca,16'h00de,16'h00af,16'h01dd,16'h001f,-16'h002c,16'h003f,16'h002a,16'h0140,16'h0011,-16'h0012,-16'h0111,16'h0063,-16'h0023,16'h00b8,-16'h0012,16'h0214,16'h00b5,-16'h003d,16'h00e7,16'h009c,16'h009d,-16'h02dd,16'h0008,16'h00aa,16'h001c,16'h01cc,-16'h00c2,-16'h0139,16'h00fe,16'h00fb,-16'h0028,-16'h0048,16'h0146,16'h0049,16'h00f8,-16'h0048,16'h0000,16'h0130,-16'h00fa,-16'h00b6,16'h019f,-16'h001b,16'h0029,-16'h0163,-16'h0007,-16'h0006,16'h0124,16'h0000,16'h0109,-16'h0099,16'h002c,-16'h00b6,16'h015c,-16'h006a,-16'h0151,-16'h0044,16'h000b,-16'h018f,-16'h00d1,-16'h004e,16'h0063,-16'h00e1,-16'h00ae,-16'h052c,16'h00ea,16'h0061,16'h01f0,16'h0084,-16'h008a,-16'h0018,16'h0090,16'h0166,16'h0091,16'h0078,-16'h00ea,-16'h0006,-16'h0064,16'h00fb,16'h003f,16'h01ee,16'h006b,16'h009f,16'h010c,-16'h0001,16'h00f7,-16'h043c,16'h00a7,16'h003e,16'h0032,16'h0068,-16'h008a,-16'h00d1,16'h0186,16'h0102,-16'h004d,16'h0012,16'h00db,16'h008f,16'h0113,-16'h002c,-16'h00b7,16'h00d8,-16'h0053,-16'h0024,16'h00d8,16'h00e4,-16'h0051,-16'h0189,-16'h004e,-16'h0058,16'h0098,-16'h0028,16'h017e,-16'h009b,-16'h0021,-16'h016a,16'h00a7,-16'h0134,-16'h0293,-16'h005f,-16'h000e,-16'h0132,-16'h00f8,-16'h00b4,16'h00e4,-16'h00c2,-16'h006f,-16'h04b2,16'h0125,-16'h0047,16'h01b3,16'h0026,-16'h0013,-16'h0061,16'h0087,16'h014e,16'h0043,16'h0020,-16'h0062,16'h00a5,-16'h0039,16'h0166,-16'h000d,16'h01d4,-16'h001a,16'h00e8,16'h0078,-16'h0066,16'h00ef,-16'h058e,16'h0018,16'h0026,16'h0154,-16'h000a,-16'h0063,-16'h00b4,16'h01c9,16'h00a7,16'h0041,16'h0050,-16'h00d5,16'h00c2,16'h0081,-16'h003b,-16'h00bb,16'h0131,-16'h0061,-16'h004b,16'h00c8,16'h0176,-16'h001a,-16'h017d,-16'h0054,-16'h0106,16'h000e,-16'h000e,16'h0289,-16'h0059,-16'h0019,-16'h01d6,16'h0007,-16'h008f,-16'h020d,16'h0024,-16'h001f,-16'h00f4,-16'h00c7,-16'h00a5,16'h00f9,-16'h00a0,-16'h01a5,-16'h00df,16'h0089,-16'h00cc,16'h01ad,-16'h000d,16'h002a,16'h0013,16'h0099,16'h01d2,16'h0034,-16'h005c,-16'h005f,16'h0159,-16'h005c,16'h01a4,-16'h0097,16'h0189,16'h0021,16'h007f,16'h011b,16'h0045,16'h005e,-16'h0637,16'h0014,16'h0010,16'h0140,-16'h00e6,16'h0029,-16'h00e4,16'h0207,-16'h0005,16'h00a3,-16'h008a,-16'h0149,16'h00d2,16'h008f,-16'h00d9,-16'h00d0,16'h00b0,-16'h0013,-16'h00c8,16'h00ef,16'h0104,-16'h00a7,-16'h0195,-16'h0006,-16'h0149,-16'h001f,16'h0064,16'h0280,-16'h00cd,-16'h002e,-16'h0170,-16'h001d,-16'h00e6,16'h0087,-16'h007f,16'h0008,-16'h0131,-16'h002f,-16'h0079,16'h0162,16'h0007,-16'h0235,16'h0055,16'h0131,-16'h0084,16'h01a2,-16'h000d,-16'h0005,-16'h007f,16'h004c,16'h01e7,-16'h0024,-16'h0051,16'h0019,16'h00f2,-16'h0041,16'h0280,-16'h007f,16'h018a,-16'h00a2,16'h005c,16'h0177,16'h004e,16'h004d,-16'h044b,16'h0050,16'h0014,16'h00fe,-16'h01ac,-16'h0041,-16'h00b3,16'h0230,16'h0012,16'h00a0,-16'h0089,-16'h01f5,16'h0079,16'h0022,-16'h00da,-16'h0077,16'h0091,-16'h0015,-16'h0027,16'h00d8,16'h0094,-16'h008a,-16'h019b,-16'h005f,-16'h0159,16'h0075,16'h00ab,16'h028d,-16'h0089,-16'h0046,-16'h010f,16'h0000,-16'h00b6,16'h0123,-16'h00db,16'h0096,-16'h0112,-16'h003e,16'h0000,16'h01b3,16'h009c,-16'h01b7,16'h0108,16'h005f,-16'h008f,16'h014d,-16'h0019,-16'h002b,-16'h00a6,16'h007d,16'h01e0,16'h0045,-16'h0082,-16'h0018,16'h0008,-16'h000f,16'h02f9,-16'h0066,16'h018f,16'h001e,16'h004a,16'h006e,-16'h0008,16'h004a,-16'h02f4,-16'h0041,16'h0077,16'h009b,-16'h0281,-16'h002e,-16'h009e,16'h024e,-16'h0003,16'h0095,16'h0020,-16'h013e,16'h0136,-16'h000f,-16'h0062,-16'h00e2,16'h0032,16'h0000,16'h007b,-16'h0070,16'h0108,-16'h0025,-16'h0153,16'h0027,-16'h00d0,16'h0094,16'h0077,16'h01fa,-16'h001b,-16'h0062,-16'h00d3,16'h0039,-16'h0117,16'h0231,-16'h011f,16'h00a7,-16'h00a9,-16'h001a,-16'h0006,16'h0121,16'h0134,-16'h0097,16'h00ff,-16'h0007,-16'h00fb,16'h01ba,16'h0010,-16'h002f,-16'h00de,16'h008e,16'h017b,16'h0000,-16'h00be,-16'h005f,-16'h01a3,16'h0060,16'h0398,-16'h00a3,16'h020e,16'h0012,16'h005a,16'h00aa,-16'h0002,16'h00c9,-16'h011c,-16'h0081,16'h0049,16'h0037,-16'h0231,-16'h0093,16'h003f,16'h028d,16'h0011,16'h009e,-16'h0021,-16'h0056,16'h0149,-16'h0013,16'h001a,-16'h0023,16'h008e,16'h0029,16'h00bd,-16'h003b,16'h00c4,16'h003b,-16'h021b,16'h0019,-16'h0130,16'h000f,16'h0082,16'h01bd,-16'h0054,-16'h001c,-16'h013a,16'h001a,-16'h00c5,16'h017c,-16'h0115,16'h0085,-16'h010c,-16'h0003,16'h0080,16'h0154,16'h01be,16'h00bc,16'h00b4,-16'h003e,-16'h006e,16'h0176,-16'h003a,-16'h0045,16'h0010,-16'h0012,16'h0194,-16'h0082,-16'h013e,-16'h00b6,-16'h022b,16'h00dc,16'h039e,16'h0015,16'h0201,16'h0028,16'h0048,16'h0031,16'h0041,16'h00f2,-16'h008e,16'h0030,16'h0070,16'h005e,-16'h01e9,-16'h0033,16'h00d6,16'h01e7,16'h0010,16'h000d,-16'h0034,16'h00c9,16'h0154,-16'h0047,16'h00cd,-16'h0068,16'h0001,-16'h006e,-16'h0018,-16'h000d,16'h00c8,16'h004e,-16'h0266,-16'h0003,-16'h00a7,-16'h0008,16'h0095,16'h016f,-16'h001c,-16'h0034,-16'h0118,-16'h0086,-16'h00cb,16'h00a5,-16'h003d,16'h0139,-16'h00f7,-16'h003a,16'h0078,16'h00be,16'h029d,16'h011d,16'h00f3,-16'h001f,16'h0030,16'h01e9,16'h006b,-16'h00aa,16'h009f,-16'h009b,16'h0186,-16'h0056,-16'h00e1,-16'h0076,-16'h021a,16'h0062,16'h0310,16'h00dc,16'h0265,16'h0030,16'h005b,16'h002a,-16'h000c,16'h0028,-16'h00bb,16'h0001,-16'h000f,16'h0068,-16'h017c,16'h003b,16'h0101,16'h0214,16'h0098,16'h001f,-16'h0070,16'h0190,16'h01d4,-16'h0028,16'h003e,16'h0008,16'h0003,-16'h001d,16'h0043,16'h002d,16'h009a,16'h0175,-16'h0261,16'h0002,-16'h00bc,16'h001a,16'h008d,16'h009f,16'h003f,-16'h0032,-16'h002b,-16'h00f0,-16'h00fa,-16'h01c4,16'h00f9,16'h015e,16'h000b,-16'h0001,16'h004f,16'h00b7,16'h024c,16'h014f,16'h0133,16'h0079,16'h006d,16'h018d,16'h0084,16'h000c,16'h005e,-16'h0060,16'h00e4,-16'h006d,-16'h008c,-16'h010d,-16'h00ce,-16'h0093,16'h0316,16'h0090,16'h024f,16'h00fe,16'h002e,16'h0053,16'h0019,16'h0008,-16'h004c,-16'h0019,-16'h0070,16'h009f,-16'h00e4,16'h00b4,16'h00ac,16'h01d7,16'h0050,16'h0030,-16'h016e,16'h014c,16'h0225,-16'h00cb,-16'h0017,-16'h0050,16'h0002,-16'h0078,16'h006c,16'h0096,16'h00a4,16'h019e,-16'h0296,-16'h0006,16'h0004,16'h00eb,16'h0066,16'h0005,16'h0061,-16'h001b,16'h001c,-16'h006a,-16'h007a,-16'h0256,16'h0112,16'h020c,16'h0055,-16'h0024,16'h0018,16'h00cb,16'h01af,16'h0185,16'h0111,16'h0033,-16'h0022,16'h01a3,16'h004c,-16'h006d,-16'h0110,-16'h000a,16'h0018,16'h0028,-16'h005a,-16'h0043,16'h00d6,-16'h0248,16'h0293,16'h0110,16'h01be,16'h0152,16'h006a,16'h002b,16'h0026,16'h0000,-16'h0060,-16'h0034,16'h001d,16'h0147,-16'h0103,16'h00e3,16'h003c,16'h0162,16'h0000,16'h008c,-16'h00fb,16'h010b,16'h0221,-16'h006f,16'h0047,-16'h00ad,16'h0016,-16'h001e,16'h0076,16'h007b,16'h001b,16'h015c,-16'h0278,16'h0064,-16'h003c,16'h00f6,16'h0099,-16'h00f0,-16'h0024,-16'h0043,16'h01bd,-16'h008a,16'h0030,-16'h0197,16'h011d,16'h01eb,16'h0041,16'h000b,-16'h006a,16'h0076,16'h0076,16'h012c,16'h0126,16'h003a,-16'h00d7,16'h0198,16'h00a8,-16'h009e,-16'h0282,16'h001e,-16'h00bb,16'h005f,-16'h0040,16'h004a,16'h006b,-16'h016f,16'h021b,16'h016b,16'h023e,16'h0069,16'h0075,-16'h0082,16'h0078,16'h0128,16'h000a,16'h000b,-16'h0004,16'h0167,-16'h012d,16'h00f6,16'h0057,16'h00fe,16'h005e,16'h00d1,-16'h011d,-16'h0002,16'h015f,-16'h003e,16'h004e,-16'h00ac,-16'h000d,-16'h0044,-16'h007d,16'h00a3,-16'h0026,16'h017b,-16'h0245,16'h000b,16'h0041,16'h0077,16'h00c3,-16'h00b3,-16'h0029,16'h001f,16'h01db,16'h0068,16'h008d,-16'h004b,16'h01cb,16'h0258,16'h0026,16'h009d,-16'h004f,16'h00b1,-16'h020d,16'h014b,16'h00a4,16'h002a,-16'h00e2,16'h00d0,16'h00c0,-16'h003a,-16'h0246,16'h0042,-16'h00b2,16'h0054,-16'h0070,16'h005d,16'h0026,16'h003a,16'h021f,16'h0180,16'h019b,16'h0009,16'h00ad,-16'h0087,16'h00c5,16'h0161,16'h00a3,16'h0006,-16'h0056,16'h01c4,-16'h00d8,16'h0184,16'h0074,16'h0148,16'h004d,16'h007f,-16'h00a0,16'h0015,16'h013f,16'h0032,16'h00bf,-16'h0082,16'h002d,-16'h005f,16'h000f,16'h0079,-16'h0082,16'h00ed,-16'h01fd,-16'h001c,16'h003f,-16'h0018,16'h0062,-16'h00fd,16'h000d,-16'h0032,16'h01c9,16'h0072,16'h0060,-16'h006a,16'h0122,16'h020f,-16'h0077,16'h0059,-16'h0016,16'h0135,-16'h05d1,16'h00dc,16'h0078,-16'h0046,-16'h0091,16'h0041,16'h00b7,-16'h004d,-16'h0161,16'h001b,-16'h00fd,16'h0011,-16'h00ac,16'h0052,-16'h0035,16'h015b,16'h023f,-16'h0002,16'h0192,-16'h00c3,16'h003e,-16'h00a1,16'h00f9,16'h00ca,16'h00e8,-16'h0089,-16'h003b,16'h00cc,-16'h0026,16'h011b,16'h0032,16'h00f1,16'h0088,16'h0029,-16'h00b9,-16'h000f,16'h016c,16'h0038,16'h00fd,-16'h0067,16'h006a,-16'h0078,16'h0039,-16'h000a,-16'h011d,16'h0115,-16'h01c8,-16'h0076,-16'h0025,-16'h0087,16'h008d,-16'h0117,-16'h0002,-16'h00d1,16'h0176,16'h0033,16'h00a5,-16'h0015,16'h0038,16'h01d7,-16'h00dd,-16'h003d,-16'h0029,16'h00f6,-16'h0882,16'h0074,-16'h0023,16'h002b,-16'h00ba,16'h005b,16'h0024,-16'h000a,16'h0002,-16'h0008,-16'h01e9,16'h0050,-16'h0031,16'h00e8,-16'h00e3,16'h019a,16'h0219,-16'h020e,16'h01a7,-16'h010c,-16'h001c,-16'h0009,16'h00bd,-16'h00d3,16'h00ad,16'h0022,-16'h0053,16'h007e,-16'h0057,16'h0097,16'h0063,16'h00a1,16'h0078,16'h0075,16'h009c,-16'h009c,16'h0102,16'h001b,16'h0089,-16'h0045,16'h00b7,-16'h002b,16'h012b,-16'h003d,-16'h01d1,16'h0148,-16'h0164,-16'h0053,16'h001c,-16'h001b,16'h0082,-16'h0151,16'h0030,-16'h005a,16'h0159,16'h00b5,16'h00f1,-16'h0017,-16'h004b,16'h012f,-16'h0138,16'h000e,-16'h000c,16'h010c,-16'h06a8,-16'h006f,-16'h0079,16'h00e9,-16'h001b,16'h006e,16'h00a6,-16'h0057,16'h0130,-16'h0047,-16'h0304,16'h0025,16'h006a,16'h0109,-16'h0075,16'h00dd,16'h0221,-16'h0265,16'h01ab,-16'h00cb,16'h0000,16'h012b,16'h00ab,-16'h03eb,16'h00fd,16'h001f,-16'h0012,16'h0080,-16'h0069,16'h001d,16'h0072,16'h0097,16'h0094,16'h00f1,16'h0106,-16'h00ae,16'h0190,-16'h0006,16'h00d4,-16'h0048,16'h00e4,-16'h002c,16'h0155,16'h0000,-16'h023f,16'h0133,-16'h0190,-16'h0063,-16'h001c,16'h00a8,16'h0056,-16'h021e,-16'h0037,-16'h004e,16'h0035,-16'h000d,16'h00b7,-16'h0026,-16'h02ab,16'h0174,-16'h0294,-16'h002e,-16'h0051,16'h00b4,-16'h031b,-16'h00b4,-16'h0071,16'h00b2,16'h0005,16'h003c,16'h0183,-16'h0105,16'h01b5,16'h003d,-16'h0387,-16'h0115,16'h00e7,16'h0109,16'h001f,-16'h0072,16'h0180,-16'h0140,16'h01ef,-16'h013b,16'h004f,16'h017d,16'h0025,-16'h05ce,16'h0146,16'h0007,-16'h0139,16'h00f8,-16'h0071,16'h0058,16'h0014,16'h00b9,16'h012b,16'h00c6,16'h0145,-16'h00d5,16'h019b,16'h0025,16'h00d9,16'h0007,16'h008b,16'h0036,16'h014e,16'h00d4,-16'h0221,16'h01a3,-16'h0185,16'h0015,16'h0031,16'h006b,16'h00e9,-16'h028b,16'h003b,16'h0026,-16'h0004,16'h0012,16'h00a1,-16'h0044,-16'h04f8,16'h013e,-16'h025b,-16'h0037,-16'h003f,16'h00be,-16'h01ab,-16'h007c,-16'h0082,16'h0093,16'h0019,-16'h0014,16'h01f5,-16'h0104,16'h00fd,-16'h006f,-16'h02c3,-16'h00b1,16'h0006,16'h009f,16'h0000,-16'h0147,16'h01a2,16'h007b,16'h0144,-16'h00cb,16'h00d7,16'h01a0,-16'h000b,-16'h06a7,16'h0169,16'h005a,-16'h00bb,16'h003b,16'h00ee,-16'h0010,-16'h0079,16'h0020,16'h0107,16'h005a,16'h0170,-16'h007d,16'h01da,16'h005a,16'h016f,16'h008a,16'h005f,16'h0085,16'h01a0,16'h00e8,-16'h01d7,16'h016e,-16'h01f2,-16'h006e,-16'h0027,16'h00c9,16'h0142,-16'h0285,16'h001a,16'h006a,-16'h00b1,16'h00a9,16'h00e3,-16'h005e,-16'h042d,16'h0120,-16'h0091,-16'h002c,-16'h0067,16'h00f8,-16'h00c9,-16'h0066,16'h0024,16'h0040,-16'h004a,-16'h004f,16'h01da,-16'h011d,-16'h0031,-16'h0083,-16'h0281,-16'h0124,-16'h00ad,16'h00c0,16'h0089,-16'h01e6,16'h0149,16'h02f2,16'h00d5,-16'h010e,16'h015e,16'h0177,16'h0064,-16'h0630,16'h00b9,16'h003b,-16'h000f,16'h00ff,16'h009a,16'h00a6,-16'h00e0,16'h0050,16'h0123,-16'h00ad,16'h0152,-16'h00f4,16'h01e0,-16'h00d6,16'h0130,16'h0139,16'h0062,16'h0084,16'h014a,16'h00eb,-16'h01c5,16'h0103,-16'h015e,-16'h000c,-16'h0022,16'h00bb,16'h00c4,-16'h02a2,16'h004e,16'h0045,-16'h0120,16'h00df,-16'h0006,-16'h0045,-16'h02cc,16'h0141,-16'h0056,16'h004f,-16'h005b,16'h00c3,-16'h00eb,-16'h004a,16'h0026,16'h0024,-16'h0021,-16'h0063,16'h0100,-16'h0062,-16'h014f,-16'h00d0,-16'h019e,-16'h00f8,-16'h0204,16'h0090,16'h004b,-16'h00ea,16'h01ec,16'h02c6,16'h0065,-16'h008c,16'h0120,16'h01b1,16'h008b,-16'h0416,16'h00af,-16'h001b,16'h001a,16'h00eb,16'h009f,16'h011c,-16'h00cb,16'h001a,16'h00f1,-16'h0263,16'h0246,-16'h00fc,16'h0207,-16'h0058,16'h0139,16'h01a7,16'h0064,-16'h000d,16'h0029,16'h0073,-16'h0212,16'h009d,-16'h00ae,-16'h000b,-16'h0047,16'h012c,16'h00f4,-16'h0231,16'h0085,16'h0106,-16'h01d8,16'h015c,-16'h0034,-16'h0075,16'h004b,16'h0120,16'h0097,16'h0034,-16'h0023,16'h0097,-16'h0066,-16'h009c,16'h004e,16'h006f,-16'h0050,-16'h00a8,16'h0001,-16'h00d4,-16'h018d,-16'h013c,-16'h00ef,-16'h0057,-16'h032f,16'h006a,-16'h00e8,16'h006e,16'h0199,16'h0316,16'h0089,-16'h007b,16'h015e,16'h0208,16'h0076,-16'h02c9,16'h0068,-16'h0002,16'h00b6,16'h0138,16'h0108,16'h010a,-16'h0062,16'h0041,16'h0052,-16'h02cb,16'h0198,-16'h007f,16'h01ae,-16'h0048,-16'h00a6,16'h00fd,-16'h00a2,-16'h0015,16'h0018,16'h00c3,-16'h01cb,16'h0004,-16'h00a2,-16'h0077,-16'h00c9,16'h0130,16'h0150,-16'h023e,16'h0048,16'h00b8,-16'h0343,16'h0144,-16'h0068,-16'h0033,16'h0238,16'h00d1,16'h017b,-16'h004a,-16'h0033,16'h00f5,-16'h00b3,-16'h00af,-16'h003d,16'h003e,-16'h008c,16'h0038,16'h00ac,-16'h00e4,-16'h01aa,-16'h003b,-16'h00b6,-16'h0031,-16'h02cc,16'h00dd,-16'h00bd,16'h0071,16'h029a,16'h01c8,16'h0011,-16'h00ce,16'h016c,16'h0238,16'h008c,-16'h0224,16'h0096,16'h0023,16'h00ad,16'h0126,16'h017b,16'h0178,-16'h00b9,-16'h0096,-16'h0029,-16'h0278,16'h01c9,-16'h00a2,16'h0193,-16'h002e,-16'h01c6,16'h012e,-16'h00a0,-16'h0008,-16'h0041,16'h00d2,-16'h0156,-16'h0098,-16'h007c,16'h000e,-16'h00d0,16'h0173,16'h0199,-16'h0195,16'h0073,16'h0023,-16'h04c5,16'h0138,-16'h003d,-16'h0058,16'h0259,16'h00cb,16'h016c,16'h002f,-16'h0048,16'h010c,-16'h007c,-16'h0080,16'h0042,-16'h0096,-16'h006c,16'h013b,16'h00c6,-16'h00d3,-16'h01ab,16'h002f,-16'h00a3,16'h0025,-16'h021a,16'h005d,-16'h009f,16'h0075,16'h0344,16'h0021,16'h00bf,-16'h0095,16'h0191,16'h0221,16'h0095,-16'h0128,16'h00b0,16'h002b,-16'h000c,16'h019b,16'h0084,16'h018b,-16'h0129,-16'h00e0,-16'h0065,-16'h01cb,16'h01a6,16'h0032,16'h019d,-16'h005c,-16'h023a,16'h0223,-16'h0045,-16'h008d,16'h0020,16'h0163,-16'h010d,-16'h0187,-16'h00b5,-16'h0003,-16'h0049,16'h003d,16'h01e3,-16'h0114,16'h0121,16'h00bc,16'h0062,16'h00ac,-16'h008f,-16'h0042,16'h00d2,16'h015e,-16'h00af,-16'h00b1,-16'h008c,-16'h000d,-16'h005b,16'h000f,16'h0289,16'h00a5,16'h0002,16'h0232,16'h00d2,-16'h00dd,16'h0012,16'h00b0,-16'h00b7,-16'h0021,-16'h0005,-16'h009d,16'h0034,-16'h0021,-16'h004e,16'h0141,16'h0112,16'h011c,-16'h00af,16'h0023,-16'h002d,16'h011a,-16'h00f4,-16'h003d,16'h00be,16'h0035,16'h0070,-16'h0117,-16'h0005,-16'h00df,16'h0044,16'h0001,16'h0110,16'h00d4,16'h0132,16'h0078,-16'h0079,-16'h0030,16'h00ea,16'h005a,16'h006a,16'h01b6,-16'h018a,-16'h0100,-16'h00a2,16'h0060,16'h002e,16'h0078,16'h00ff,-16'h011a,16'h0091,16'h012b,-16'h0089,16'h0092,-16'h0014,-16'h0005,-16'h003e,16'h00dc,-16'h0096,-16'h0085,-16'h00ef,-16'h0037,-16'h003b,-16'h004d,16'h014f,16'h009c,-16'h0062,16'h0245,16'h0073,-16'h00cd,16'h0042,16'h0051,-16'h00df,-16'h0008,-16'h002a,-16'h000b,16'h0010,-16'h00a1,-16'h0047,16'h0027,16'h0115,16'h0085,-16'h0121,-16'h0085,-16'h0048,16'h00e4,-16'h01ff,-16'h0070,16'h008c,16'h0070,16'h0171,16'h0046,-16'h00d4,-16'h00e5,16'h00af,16'h006b,16'h00a4,16'h00bc,16'h008b,16'h0090,-16'h0056,-16'h0046,16'h00fa,16'h0070,-16'h00a7,16'h013c,-16'h023b,-16'h006c,-16'h0156,16'h0122,16'h0009,16'h00ad,16'h00a8,-16'h024d,-16'h000a,16'h01a7,-16'h007e,16'h0098,-16'h0075,16'h0152,-16'h0086,16'h0106,-16'h0121,-16'h00b9,-16'h00c8,16'h0055,-16'h0033,-16'h0113,16'h00b8,16'h005d,-16'h00b2,16'h01e6,-16'h001d,-16'h001c,-16'h0070,16'h003c,-16'h0066,16'h000b,16'h0026,-16'h0069,-16'h004c,-16'h00f8,-16'h0078,-16'h0036,16'h00de,16'h00ae,-16'h01b1,16'h0032,16'h005e,16'h00f0,-16'h0285,-16'h0085,16'h0095,-16'h003a,16'h017a,16'h00f0,-16'h011e,-16'h00f7,16'h0077,16'h0001,16'h0042,16'h013e,16'h00a1,16'h009a,16'h0000,-16'h0079,16'h011d,-16'h005f,-16'h00c7,16'h0091,-16'h0239,-16'h005a,-16'h01ac,16'h0105,-16'h005c,16'h0074,16'h0078,-16'h0237,-16'h0076,16'h013f,-16'h0036,16'h0110,-16'h002d,16'h0165,-16'h0099,16'h0050,-16'h0174,-16'h0040,-16'h008f,-16'h0032,-16'h0040,-16'h01b6,-16'h0008,16'h0012,-16'h006e,16'h0217,16'h006b,-16'h0035,-16'h0002,16'h005d,-16'h004b,-16'h0004,-16'h00b0,-16'h001a,-16'h008c,-16'h002d,-16'h001e,16'h001f,16'h01a0,16'h0184,-16'h01df,16'h001f,-16'h0006,16'h00cc,-16'h0301,-16'h0085,16'h0080,16'h008f,16'h020c,16'h009d,-16'h016b,-16'h0093,16'h0045,16'h0016,16'h00f2,16'h016f,16'h0081,16'h00d2,-16'h0026,-16'h0036,16'h0158,-16'h0074,-16'h00e1,16'h008f,-16'h00f9,-16'h005f,-16'h0248,16'h0127,-16'h0065,16'h00d8,16'h008e,-16'h00da,-16'h004b,16'h00dc,-16'h0070,16'h014b,-16'h009c,16'h0061,-16'h00e5,16'h0051,-16'h0264,-16'h0071,-16'h00d5,16'h0052,-16'h007b,-16'h01a4,-16'h015c,16'h00a7,-16'h003f,16'h01df,16'h0017,-16'h008c,-16'h000e,16'h0074,16'h004c,-16'h0081,-16'h0091,16'h0008,-16'h0064,-16'h009a,16'h0025,-16'h0059,16'h013d,16'h00fe,-16'h0128,16'h0000,-16'h000b,16'h00c2,-16'h02ed,-16'h003d,16'h0099,16'h0139,16'h0207,16'h0034,-16'h01d5,-16'h009a,16'h001f,-16'h0026,16'h00e9,16'h015e,16'h0102,16'h0186,-16'h0035,-16'h001c,16'h0104,-16'h0089,-16'h0123,16'h00d4,-16'h0056,-16'h0057,-16'h0253,16'h0170,-16'h005a,16'h0103,16'h008e,-16'h002f,-16'h00c8,-16'h0027,16'h0028,16'h00d0,-16'h005d,-16'h0039,-16'h00c2,16'h0083,-16'h02be,-16'h00a4,-16'h00eb,16'h0047,-16'h00ed,-16'h011f,-16'h0304,16'h012f,16'h006f,16'h030e,16'h007f,-16'h00a8,16'h0010,16'h0038,16'h0109,-16'h0004,-16'h001d,-16'h00c3,16'h005b,-16'h0077,-16'h0040,16'h0043,16'h0135,16'h009c,16'h0022,16'h0040,16'h0048,16'h0102,-16'h03b2,-16'h0016,16'h0075,16'h014e,16'h01bd,16'h0071,-16'h0159,-16'h001f,16'h0115,-16'h004a,16'h00ca,16'h009a,16'h00cc,16'h014d,-16'h00c7,-16'h0027,16'h00dc,-16'h0097,-16'h013a,16'h00e8,16'h00b7,-16'h007d,-16'h01a2,16'h0109,16'h0033,16'h00e0,16'h0008,16'h014a,-16'h00c6,-16'h0021,-16'h0096,16'h00f8,-16'h004a,-16'h0297,-16'h0065,16'h00cb,-16'h0305,-16'h006f,-16'h0170,16'h00af,-16'h007e,-16'h00a2,-16'h044c,16'h00fa,16'h0019,16'h0295,16'h0092,-16'h007e,-16'h0090,16'h0148,16'h00e7,16'h0031,-16'h0076,-16'h008b,16'h006d,-16'h00e3,16'h0029,16'h0076,16'h00f6,16'h0009,16'h00bb,16'h00a6,16'h0079,16'h0143,-16'h0515,16'h004b,16'h00f3,16'h0195,16'h010f,16'h000e,-16'h012b,16'h00cd,16'h014f,-16'h0074,16'h00c3,-16'h0090,16'h00c1,16'h0092,-16'h0066,16'h000d,16'h011b,-16'h008b,-16'h00f2,16'h00bb,16'h0130,-16'h00bd,-16'h013d,16'h00f9,-16'h0017,16'h00b8,16'h0071,16'h01f8,-16'h0094,-16'h0051,-16'h0172,16'h0098,-16'h0077,-16'h036e,-16'h000d,-16'h0011,-16'h0222,-16'h0104,-16'h013b,16'h00e4,-16'h00b5,-16'h0137,-16'h0291,16'h00b6,16'h000f,16'h029a,16'h00cc,-16'h003c,-16'h0025,16'h0164,16'h00f9,16'h0012,16'h0039,-16'h00a8,16'h015b,-16'h0094,16'h0023,16'h005a,16'h00d4,-16'h00d6,16'h00c6,16'h00a3,16'h00cc,16'h00a0,-16'h0582,16'h000b,16'h0039,16'h024a,16'h0014,16'h0024,-16'h010b,16'h01a1,16'h00eb,16'h0024,16'h00e3,-16'h0132,16'h007e,16'h0057,-16'h009d,-16'h001b,16'h00cd,-16'h0007,-16'h00cb,16'h0018,16'h0139,-16'h0110,-16'h009a,16'h0079,-16'h00c5,16'h0094,16'h005f,16'h01bf,-16'h009e,-16'h00b6,-16'h0206,16'h0024,-16'h0086,-16'h0169,-16'h0085,16'h000b,-16'h020d,-16'h00a0,-16'h0112,16'h00f0,16'h0014,-16'h0242,16'h0010,16'h009a,-16'h005b,16'h025c,-16'h0072,16'h0040,-16'h001e,16'h00a7,16'h0175,16'h0012,-16'h002b,-16'h000c,16'h01eb,-16'h0053,16'h001a,-16'h0017,16'h0073,-16'h00cf,16'h0042,16'h006e,16'h0035,16'h0094,-16'h04c4,-16'h003f,16'h0061,16'h0233,-16'h00dc,16'h0060,-16'h00f6,16'h0261,16'h0005,-16'h0017,16'h00e5,-16'h0164,16'h0048,-16'h0040,-16'h0064,-16'h0007,16'h00b5,-16'h0055,-16'h0024,16'h0060,16'h00ae,-16'h0115,-16'h004c,16'h006e,-16'h00bb,16'h0029,16'h00d6,16'h01d9,-16'h00e9,-16'h007d,-16'h0201,16'h0026,-16'h00d2,16'h00f7,-16'h00a9,16'h009c,-16'h0204,-16'h0057,-16'h00fb,16'h019b,16'h0013,-16'h01cc,16'h00ec,-16'h001d,-16'h0106,16'h01c6,16'h0001,-16'h000a,-16'h00a2,16'h0029,16'h021f,16'h004b,16'h0005,-16'h003a,16'h00e2,-16'h005d,16'h00fb,-16'h0080,16'h0073,-16'h00b7,16'h0087,16'h00fd,16'h0022,16'h0076,-16'h02ea,-16'h0076,16'h0098,16'h01f8,-16'h0203,16'h002a,-16'h0117,16'h02d8,-16'h0094,16'h003c,16'h00c7,-16'h0140,16'h0082,-16'h0074,-16'h00cf,-16'h0015,16'h0082,-16'h0040,16'h002c,16'h0035,16'h00cd,-16'h00e1,16'h0022,16'h0042,-16'h0074,16'h0093,16'h00ea,16'h0170,-16'h00ae,-16'h00b2,-16'h014f,16'h0038,-16'h00f3,16'h024a,-16'h00ba,16'h00de,-16'h00a7,-16'h0040,-16'h00b0,16'h012e,16'h00af,-16'h00e7,16'h00d8,16'h003e,-16'h00e0,16'h018d,16'h001c,-16'h0030,-16'h007b,16'h0052,16'h01f8,-16'h0038,-16'h0023,-16'h0056,-16'h0092,-16'h004c,16'h01c9,-16'h004f,16'h00a0,-16'h0099,16'h00ba,16'h00a7,-16'h004d,16'h0110,-16'h01c9,-16'h004b,16'h005c,16'h0174,-16'h0282,16'h000d,-16'h0107,16'h0342,-16'h002a,16'h00a0,16'h0069,-16'h0040,16'h00ba,-16'h007f,-16'h0020,-16'h003b,16'h00f6,-16'h0067,16'h00b8,16'h002c,16'h00d2,-16'h001d,-16'h0021,16'h0065,-16'h0054,16'h0068,16'h00cc,16'h0142,-16'h00ce,-16'h00bd,-16'h00ea,16'h002a,-16'h0136,16'h024e,-16'h0119,16'h00cc,-16'h0054,-16'h0035,-16'h0039,16'h0156,16'h017d,-16'h00ca,16'h0110,16'h0003,-16'h0049,16'h01f0,-16'h0029,16'h000c,-16'h0076,16'h0029,16'h015c,-16'h00f8,-16'h008b,-16'h00f5,-16'h021e,16'h00ce,16'h02d5,-16'h0085,16'h0082,-16'h0070,16'h0083,16'h0081,-16'h011a,16'h00c9,-16'h0073,-16'h0037,16'h004e,16'h017f,-16'h01eb,-16'h001c,16'h001f,16'h033d,16'h004c,16'h00cb,16'h00b1,-16'h0001,16'h00be,-16'h009d,16'h0038,-16'h001a,16'h0058,-16'h003b,16'h0065,16'h0005,16'h0024,-16'h0007,16'h000a,16'h0075,-16'h0035,16'h0042,16'h0106,16'h018d,-16'h0052,-16'h0036,-16'h0067,-16'h000b,-16'h00f7,16'h0195,-16'h00fd,16'h0162,-16'h0127,-16'h0035,16'h001a,16'h013e,16'h01c5,16'h005e,16'h0107,-16'h0054,16'h0001,16'h0213,-16'h002f,-16'h008c,16'h004c,-16'h0058,16'h01b3,-16'h00e3,-16'h010a,-16'h0124,-16'h0209,16'h019a,16'h0301,16'h004c,16'h009b,16'h0055,16'h000d,-16'h0014,-16'h0105,-16'h0032,-16'h0059,-16'h00a2,16'h005a,16'h01c8,-16'h01ad,16'h003f,16'h00d5,16'h0388,16'h008b,16'h00a8,16'h0036,16'h0144,16'h015d,-16'h00af,16'h00bb,-16'h0065,16'h005d,16'h0000,16'h0003,16'h002d,-16'h00a6,16'h00e2,-16'h0058,16'h004c,-16'h001d,16'h000c,16'h00a2,16'h017b,16'h0016,-16'h00c9,-16'h00ba,-16'h0068,-16'h00fc,-16'h005e,-16'h0030,16'h012c,-16'h0149,-16'h0027,-16'h002b,16'h010f,16'h018d,16'h0080,16'h00da,16'h0021,16'h003f,16'h021e,-16'h0062,-16'h0021,16'h009b,-16'h00ad,16'h00cc,-16'h0111,-16'h008c,-16'h00cb,-16'h013e,16'h0114,16'h0318,16'h008d,16'h0081,16'h00a2,-16'h0081,-16'h006e,-16'h00db,-16'h00b3,-16'h0099,-16'h0022,-16'h001c,16'h0147,-16'h0144,16'h0112,16'h0095,16'h0342,-16'h000c,16'h004b,-16'h0020,16'h017e,16'h0126,-16'h00af,16'h0083,-16'h0072,16'h006a,-16'h0023,16'h0087,16'h0092,-16'h01cb,16'h0078,-16'h0094,16'h0031,-16'h0047,16'h00a4,16'h0110,16'h009e,16'h0074,-16'h00ff,-16'h005d,-16'h00ca,-16'h0101,-16'h031c,16'h007f,16'h0167,-16'h0070,-16'h0009,16'h0027,16'h00de,16'h01b0,16'h0104,16'h0196,16'h002f,16'h00dd,16'h0234,16'h0032,16'h0020,16'h0053,-16'h007d,16'h001c,-16'h00d7,-16'h00a9,-16'h0059,-16'h003d,-16'h00bd,16'h02db,16'h006d,16'h0145,16'h00ed,-16'h001c,16'h001c,-16'h0028,-16'h00e5,-16'h00d0,-16'h00be,-16'h0078,16'h01b2,-16'h00f6,16'h00ec,16'h0099,16'h032e,16'h0031,-16'h004c,-16'h004b,16'h0101,16'h0162,-16'h006d,16'h00cf,-16'h0049,16'h0059,-16'h0001,16'h00f3,16'h0023,-16'h0231,16'h00d3,-16'h0141,16'h0027,16'h001b,16'h0121,16'h0107,-16'h0026,16'h0077,-16'h00f4,16'h00be,-16'h004f,-16'h00fc,-16'h0255,16'h00ea,16'h0172,16'h0047,-16'h0012,16'h002b,16'h009e,16'h00fb,16'h0119,16'h0192,-16'h0004,-16'h0022,16'h01b9,16'h0058,-16'h0064,-16'h00b2,-16'h0023,-16'h00f0,-16'h0068,-16'h0043,16'h009d,16'h008c,-16'h02c5,16'h02e1,16'h0073,16'h0124,16'h00ab,16'h009e,-16'h000d,16'h0009,-16'h0028,16'h000d,-16'h0015,-16'h00d9,16'h0190,-16'h0066,16'h012a,16'h0033,16'h0261,-16'h006c,-16'h0090,-16'h0094,16'h0102,16'h014d,-16'h0089,16'h009d,-16'h0060,16'h0007,-16'h0024,16'h0060,16'h00a9,-16'h02cb,16'h016c,-16'h0106,16'h0006,-16'h000d,16'h0173,16'h0128,-16'h00d6,16'h0067,-16'h00ed,16'h020e,-16'h0003,-16'h000d,-16'h0125,16'h00d2,16'h0188,16'h004d,-16'h000e,-16'h0045,16'h00df,-16'h0023,16'h0118,16'h013b,16'h0038,-16'h0024,16'h019b,16'h006f,-16'h0052,-16'h01ec,16'h0044,-16'h013f,16'h0098,-16'h0065,16'h0037,16'h00f1,-16'h01c2,16'h02e7,16'h0123,16'h0121,16'h0011,16'h0036,-16'h0078,-16'h0070,16'h0077,16'h0002,16'h0006,-16'h00eb,16'h025e,16'h001e,16'h00ca,16'h00a3,16'h0251,-16'h0031,-16'h004c,-16'h00ad,16'h003b,16'h0131,-16'h0081,16'h0065,-16'h007f,-16'h000d,-16'h008d,-16'h0059,16'h0087,-16'h0348,16'h00fb,-16'h0094,-16'h0050,16'h0049,16'h0127,16'h0110,-16'h00c2,16'h0082,-16'h00bd,16'h01ea,-16'h000e,-16'h006c,-16'h007a,16'h00a3,16'h0159,-16'h0006,16'h000d,-16'h0035,16'h008c,-16'h01c6,16'h0143,16'h002b,16'h009e,-16'h004b,16'h0097,16'h00e8,-16'h0047,-16'h024b,16'h00b9,-16'h014f,16'h00b4,-16'h002e,16'h006d,16'h0004,16'h007b,16'h02ce,16'h0104,16'h00ed,-16'h0080,16'h0034,-16'h00b2,-16'h0008,16'h0118,16'h00b9,16'h0016,-16'h00bf,16'h019f,16'h00d1,16'h00bf,16'h0045,16'h021e,16'h0019,16'h0059,-16'h00d6,-16'h0085,16'h015a,-16'h0009,16'h0086,-16'h0043,-16'h0003,-16'h0098,-16'h003f,16'h009c,-16'h0409,16'h008f,-16'h0028,-16'h0001,16'h0031,16'h0032,16'h00d4,-16'h00b0,16'h00a0,-16'h007b,16'h01b5,16'h0040,-16'h0047,-16'h002a,16'h00d8,16'h01ac,16'h0093,16'h00a0,-16'h0017,16'h00c5,-16'h0539,16'h00ec,-16'h0027,16'h0057,-16'h0023,16'h00b7,16'h00bf,-16'h0032,-16'h01e8,-16'h0001,-16'h0129,16'h0099,-16'h0098,16'h003d,-16'h000c,16'h01a3,16'h02fa,-16'h0053,16'h005c,-16'h00f7,16'h002f,-16'h00af,16'h0010,16'h0151,16'h0056,16'h002f,-16'h00a8,16'h016f,16'h00b1,16'h009f,-16'h0015,16'h016e,-16'h0004,16'h0099,-16'h007d,-16'h01aa,16'h020c,16'h007b,16'h0099,-16'h0036,16'h003f,-16'h00a0,-16'h0026,-16'h000e,-16'h0429,16'h00ae,-16'h0001,16'h0052,-16'h0078,16'h0006,16'h0129,-16'h00a9,16'h0073,-16'h00a2,16'h0131,16'h0110,-16'h0025,16'h0075,-16'h0027,16'h0121,16'h001b,16'h0044,-16'h007f,16'h0083,-16'h0781,16'h007f,-16'h001c,16'h0047,-16'h0021,16'h00ca,16'h00cc,-16'h0044,-16'h00b4,-16'h0043,-16'h0200,16'h0095,-16'h0078,16'h0089,-16'h005c,16'h0157,16'h030e,-16'h020c,16'h0044,-16'h0173,-16'h002c,-16'h00b7,16'h001c,16'h0039,16'h0096,16'h0097,-16'h00aa,16'h013b,16'h0089,16'h006c,16'h0036,16'h01b4,-16'h002e,16'h0095,16'h001c,-16'h0148,16'h021c,16'h006a,16'h006c,-16'h001d,16'h002b,-16'h00dc,16'h000b,-16'h003d,-16'h04e2,16'h00ac,16'h0026,16'h000c,16'h0005,-16'h0029,16'h00c6,-16'h0091,16'h0010,-16'h004a,16'h0098,16'h0064,16'h0023,16'h0021,-16'h012a,16'h0135,-16'h012d,-16'h0026,-16'h0078,16'h00be,-16'h0643,-16'h000c,-16'h0094,16'h000c,-16'h0075,16'h0124,16'h009e,-16'h0023,16'h016c,16'h0029,-16'h02d4,-16'h0053,-16'h005d,16'h017c,-16'h0008,16'h0127,16'h022a,-16'h02c4,16'h0026,-16'h019b,-16'h0018,-16'h0059,16'h000b,-16'h015d,16'h0048,16'h00b6,-16'h00e0,16'h0159,-16'h00a7,16'h0019,16'h00b9,16'h0179,16'h0105,16'h0103,16'h0106,-16'h00c5,16'h01f0,16'h006c,16'h0081,16'h0009,16'h00d3,-16'h00b1,16'h00d7,16'h0064,-16'h04d4,16'h00d2,16'h004a,16'h003d,-16'h003d,16'h0081,16'h0164,-16'h00dd,-16'h000d,-16'h0021,16'h0054,16'h0066,16'h0093,16'h0009,-16'h02b4,16'h01a8,-16'h0253,-16'h009e,-16'h0021,16'h005d,-16'h0364,-16'h00d1,-16'h00c3,-16'h0043,16'h0027,16'h0138,16'h00b3,-16'h002a,16'h020c,-16'h004b,-16'h0376,-16'h0172,16'h009d,16'h016e,16'h0009,-16'h0021,16'h0245,-16'h00fc,16'h0000,-16'h0190,16'h0012,16'h00f7,16'h0047,-16'h02e6,16'h002b,16'h0143,-16'h01c5,16'h00d9,-16'h0086,-16'h001b,-16'h0014,16'h0122,16'h0068,16'h00da,16'h0149,-16'h00ae,16'h0158,16'h0003,16'h015b,-16'h0011,16'h00e7,-16'h0052,16'h0164,16'h00da,-16'h04d6,16'h010d,16'h0023,16'h0031,-16'h005b,16'h00e2,16'h0188,-16'h0189,16'h0056,16'h005a,-16'h008b,16'h000c,16'h00c3,-16'h005b,-16'h0598,16'h0178,-16'h0281,-16'h0075,-16'h0057,16'h0043,-16'h01b1,-16'h003e,-16'h0067,-16'h002e,16'h0059,16'h00d4,16'h0166,-16'h0019,16'h01aa,-16'h006f,-16'h023c,-16'h0209,16'h0064,16'h0159,16'h0063,-16'h011e,16'h01df,16'h006d,16'h0062,-16'h01ce,16'h00b1,16'h01b2,16'h00a2,-16'h04e0,-16'h000d,16'h00f2,-16'h0125,16'h0135,16'h000b,-16'h0003,-16'h005d,16'h00c4,16'h0051,16'h0103,16'h0177,-16'h0082,16'h01eb,-16'h004c,16'h01fb,16'h0078,16'h003b,16'h0005,16'h0108,16'h00df,-16'h0432,16'h0156,-16'h0014,16'h001e,16'h0012,16'h00e5,16'h018f,-16'h034d,16'h0087,16'h00c6,-16'h00b1,16'h003d,16'h00c6,-16'h0005,-16'h0522,16'h00d1,-16'h01d0,-16'h0096,-16'h00e4,16'h00d8,-16'h0181,-16'h0045,-16'h005a,16'h0059,-16'h000f,16'h0034,16'h014b,-16'h009b,16'h002f,-16'h0032,-16'h01d3,-16'h010a,-16'h004a,16'h0127,16'h001d,-16'h0167,16'h0249,16'h028f,16'h0052,-16'h0147,16'h00d0,16'h010c,16'h00a9,-16'h0635,-16'h0039,16'h00bc,-16'h0086,16'h0121,16'h002e,16'h0058,-16'h00e9,16'h0044,16'h00ce,-16'h008d,16'h01aa,-16'h00c0,16'h024f,-16'h00e2,16'h01e4,16'h0091,16'h0019,16'h0016,16'h00cd,16'h00e6,-16'h03ee,16'h00b2,-16'h004d,16'h004d,-16'h0073,16'h0087,16'h019f,-16'h0350,16'h00c9,16'h010b,-16'h0127,16'h008c,-16'h000e,16'h0085,-16'h0332,16'h008c,-16'h0085,-16'h0050,-16'h0092,16'h00e8,-16'h0119,-16'h0008,-16'h004d,16'h000b,16'h0020,-16'h0010,16'h00b9,-16'h0093,-16'h0137,-16'h0051,-16'h00f5,-16'h00e0,-16'h01e2,16'h0094,-16'h009f,-16'h00ac,16'h025e,16'h0319,16'h0072,-16'h01cf,16'h014f,16'h0175,16'h00c6,-16'h054b,-16'h006b,-16'h000d,-16'h003d,16'h013d,16'h00b6,16'h003d,-16'h00d5,16'h0009,16'h00a1,-16'h01be,16'h020e,-16'h00bc,16'h0259,-16'h0091,16'h0088,16'h00f5,-16'h0010,16'h0033,16'h00ae,16'h0049,-16'h034e,-16'h005c,-16'h00a4,-16'h000f,-16'h00ce,16'h00f3,16'h01ca,-16'h02e0,16'h010f,16'h0153,-16'h01a9,16'h0144,-16'h00e0,-16'h002f,-16'h002b,16'h0091,16'h008e,-16'h007d,-16'h00b0,16'h0113,-16'h0094,-16'h0069,-16'h00ec,16'h00b5,-16'h00aa,-16'h0008,16'h0023,-16'h0027,-16'h014d,-16'h0111,-16'h0089,-16'h0071,-16'h0331,16'h0043,-16'h009a,16'h005f,16'h0233,16'h0336,16'h0072,-16'h0147,16'h0113,16'h0214,16'h00da,-16'h0306,-16'h010c,-16'h004a,16'h005f,16'h013f,16'h00ea,16'h0037,-16'h002e,-16'h002a,16'h0006,-16'h01d3,16'h0234,-16'h0037,16'h01c6,-16'h004f,-16'h0149,16'h0052,16'h002c,16'h003e,16'h001d,16'h002b,-16'h02b7,-16'h0047,-16'h0176,-16'h004b,-16'h00aa,16'h0120,16'h0183,-16'h01d4,16'h00a5,16'h0127,-16'h02c4,16'h0148,-16'h0013,16'h0004,16'h019f,16'h0030,16'h0186,16'h0014,-16'h00c0,16'h011c,-16'h00dc,16'h0005,-16'h0069,16'h0088,-16'h0059,16'h00ab,16'h005d,-16'h00d4,-16'h0144,-16'h00c4,16'h0001,-16'h0079,-16'h0318,-16'h000e,-16'h00e3,16'h00c4,16'h0288,16'h021e,16'h0075,-16'h018d,16'h00af,16'h0273,16'h008e,-16'h0266,-16'h00d1,-16'h009a,16'h0122,16'h0165,16'h0117,16'h00de,-16'h00cb,-16'h00f3,-16'h006d,-16'h0180,16'h01c4,-16'h00a1,16'h019b,-16'h003b,-16'h01c5,16'h0045,-16'h0067,-16'h0005,16'h005e,16'h00d5,-16'h0261,-16'h00e0,-16'h014e,-16'h00cb,-16'h0165,16'h016d,16'h01bb,-16'h0155,16'h008e,16'h00a3,-16'h03bf,16'h0151,16'h00b1,-16'h005d,16'h02c7,16'h0014,16'h01b2,16'h0046,-16'h00f6,16'h019c,-16'h0081,16'h0000,-16'h006c,16'h0016,-16'h0134,16'h00f5,16'h0001,-16'h0086,-16'h0167,-16'h0005,-16'h002b,16'h0086,-16'h029f,16'h00c3,-16'h00d2,16'h00d6,16'h034a,16'h00e5,16'h0067,-16'h00f9,16'h014b,16'h025e,16'h0074,-16'h019e,-16'h0067,-16'h002c,16'h0097,16'h01cc,16'h006b,16'h019c,-16'h01a9,-16'h016a,-16'h008e,-16'h0161,16'h01a4,-16'h001a,16'h0193,-16'h0068,-16'h0227,16'h0205,-16'h00da,-16'h0025,-16'h0044,16'h0106,-16'h011f,-16'h00b4,-16'h00ef,16'h0007,-16'h0120,16'h000a,16'h0213,-16'h00fe,16'h008e,16'h004e,16'h0083,16'h00fa,-16'h007b,-16'h000e,16'h004d,16'h00e5,-16'h0087,-16'h00b9,-16'h003b,-16'h0023,16'h0028,16'h008d,16'h01b6,16'h0120,-16'h00b7,16'h01f5,16'h00e7,-16'h00d2,16'h0012,16'h004d,-16'h0092,-16'h004b,-16'h00c9,-16'h00c6,16'h005b,-16'h0031,-16'h00d7,16'h00e0,16'h00c4,16'h00e5,-16'h0190,16'h0043,16'h003b,16'h015b,-16'h0111,-16'h008e,16'h006b,-16'h0023,16'h009e,16'h0016,16'h0006,-16'h0157,16'h0060,-16'h0012,16'h00ca,16'h016f,16'h00d1,16'h00a8,-16'h0033,-16'h0091,16'h0054,16'h00a9,16'h005a,16'h01b3,-16'h01ec,-16'h00fc,-16'h0091,16'h00c7,-16'h00e2,16'h004f,16'h0106,-16'h0183,16'h0056,16'h0121,16'h0002,16'h00ae,-16'h0021,16'h0092,16'h0012,16'h00e3,-16'h0032,-16'h00c5,-16'h00b5,-16'h005e,16'h003c,-16'h008c,16'h0002,16'h0076,-16'h0087,16'h0207,16'h004f,-16'h0086,-16'h0037,16'h0026,-16'h012c,-16'h000f,-16'h00fc,-16'h0006,-16'h005a,-16'h00d3,-16'h00d6,16'h000d,-16'h0004,16'h0089,-16'h01d7,16'h0005,16'h00e5,16'h0131,-16'h0182,-16'h0033,16'h0067,16'h0029,16'h0110,16'h0107,-16'h00fa,-16'h010b,16'h00d9,-16'h0018,16'h0063,16'h00ee,16'h00a0,16'h0073,-16'h0013,-16'h00bc,16'h00c4,16'h0073,-16'h0006,16'h00f1,-16'h0207,-16'h0047,-16'h00fc,16'h010d,-16'h0061,16'h0029,16'h0083,-16'h01e6,-16'h0050,16'h00c9,-16'h00c4,16'h00eb,-16'h0061,16'h014d,-16'h0063,16'h010a,-16'h0114,-16'h0087,-16'h0054,16'h0019,-16'h0006,-16'h023a,-16'h001c,16'h0011,-16'h0080,16'h01fe,16'h001c,-16'h0056,-16'h0001,16'h0013,-16'h00d4,16'h000a,-16'h0079,16'h007a,16'h0000,-16'h0091,-16'h0079,16'h006b,16'h006a,16'h0137,-16'h01f1,16'h0010,16'h0076,16'h014f,-16'h01f8,-16'h00ae,16'h007f,16'h0131,16'h0116,16'h011c,-16'h00d6,-16'h00a5,16'h005e,16'h0045,16'h008c,16'h0169,16'h0009,16'h00bf,16'h0089,-16'h006f,16'h0041,-16'h0031,-16'h011c,16'h010e,-16'h00fe,-16'h00f3,-16'h0144,16'h0114,-16'h00e0,16'h006d,16'h00b0,-16'h01c3,16'h0040,16'h00ac,-16'h0089,16'h0074,16'h001d,16'h012c,-16'h0111,16'h00d9,-16'h01bc,-16'h0095,-16'h00fd,16'h0073,16'h0043,-16'h0295,-16'h0078,-16'h0039,16'h0023,16'h016e,-16'h006b,-16'h007d,-16'h0013,16'h0038,-16'h0078,16'h000b,-16'h00b8,-16'h0035,-16'h0061,-16'h0002,-16'h0035,-16'h0040,16'h00fb,16'h00fd,-16'h0175,16'h003e,16'h00ca,16'h00b1,-16'h023d,-16'h00ac,16'h0084,16'h016b,16'h0185,16'h0110,-16'h018d,-16'h00d6,-16'h000d,16'h0026,16'h00cc,16'h017c,16'h00b4,16'h0160,16'h0069,-16'h00b2,16'h0055,-16'h002f,-16'h0132,16'h00e4,-16'h00cf,-16'h006c,-16'h01d2,16'h0149,-16'h00b6,16'h0047,16'h006b,-16'h003c,16'h0031,16'h0030,-16'h00cb,16'h005c,16'h000e,16'h0066,-16'h00bf,16'h00d0,-16'h0276,-16'h0082,-16'h00b1,16'h0066,-16'h003f,-16'h01b3,-16'h0231,16'h0026,16'h0040,16'h0197,16'h009d,-16'h005e,16'h0044,16'h0037,16'h0094,-16'h000e,-16'h009c,16'h0034,-16'h0072,-16'h0061,16'h0054,16'h0005,16'h00e5,16'h00f0,-16'h00e3,-16'h0025,16'h005e,16'h0102,-16'h02c6,-16'h0043,16'h006c,16'h0153,16'h013e,16'h00c4,-16'h01c7,-16'h00c7,16'h0082,-16'h0002,16'h0116,16'h01bd,16'h0151,16'h0179,-16'h003f,-16'h0010,-16'h001f,-16'h003c,-16'h00e4,16'h00f9,16'h00a6,-16'h00a2,-16'h0130,16'h0151,-16'h0022,16'h0018,16'h0087,16'h00a9,-16'h004c,-16'h003a,-16'h001a,16'h00c7,16'h0019,-16'h00b6,-16'h00a1,16'h00cf,-16'h0221,-16'h005f,-16'h0135,16'h0084,-16'h00c3,-16'h012b,-16'h03a7,16'h0000,16'h0084,16'h0256,16'h007f,-16'h00cd,16'h002e,16'h0033,16'h007c,-16'h005a,-16'h00d2,-16'h0084,-16'h0063,-16'h00a9,16'h001a,16'h0034,16'h006d,16'h011a,16'h004e,-16'h0020,16'h002e,16'h0104,-16'h038c,-16'h0006,16'h00a3,16'h01e3,16'h01b8,16'h00db,-16'h017d,-16'h014c,16'h00f6,-16'h0045,16'h010d,16'h00e0,16'h007b,16'h00ee,16'h0017,-16'h0014,16'h0041,-16'h0036,-16'h0128,16'h00b9,16'h00d4,-16'h00ca,-16'h015e,16'h01ad,16'h0046,16'h009d,16'h002a,16'h01e2,-16'h0103,-16'h00bb,-16'h0064,16'h0041,-16'h0042,-16'h02c0,-16'h0097,16'h0096,-16'h01a2,-16'h005b,-16'h0108,16'h0028,-16'h0033,-16'h00d4,-16'h033d,16'h0086,-16'h0018,16'h02af,16'h0018,-16'h00e9,-16'h0039,16'h00b8,16'h00dc,-16'h00a2,-16'h0028,-16'h00d2,16'h00de,-16'h0066,-16'h00a0,16'h00b2,16'h005a,-16'h00b9,16'h00b6,-16'h000b,16'h0043,16'h012a,-16'h0413,16'h001a,16'h0056,16'h0242,16'h00f1,16'h0106,-16'h0108,-16'h012f,16'h00d5,-16'h0049,16'h00ed,-16'h008b,-16'h0018,16'h003a,-16'h005d,16'h0027,16'h0058,-16'h0007,-16'h00c4,16'h0086,16'h012d,-16'h0141,-16'h00df,16'h01d0,16'h00b2,16'h0022,16'h005b,16'h01a8,-16'h007d,-16'h00ae,-16'h00e6,16'h0053,-16'h0009,-16'h02c3,-16'h008d,16'h008f,-16'h01b0,-16'h0056,-16'h00f7,16'h006e,-16'h001e,-16'h0199,-16'h0066,16'h00cd,16'h001d,16'h0285,16'h0033,-16'h00a9,-16'h0081,16'h00e7,16'h012e,-16'h0095,-16'h001d,-16'h00b2,16'h0231,-16'h0170,-16'h00a1,16'h002c,-16'h002f,-16'h00ea,-16'h000c,16'h0063,16'h006d,16'h0122,-16'h03a8,16'h000f,16'h0023,16'h029c,16'h0009,16'h0124,-16'h012a,-16'h0089,16'h007a,-16'h00a7,16'h016e,-16'h0150,16'h005c,-16'h002d,-16'h0064,-16'h000f,16'h0100,-16'h00c7,-16'h00c2,16'h0000,16'h00c4,-16'h018c,-16'h0005,16'h01d7,16'h00c5,16'h0001,16'h00fe,16'h0173,-16'h00b6,-16'h00cd,-16'h009b,16'h000a,16'h001e,-16'h0010,-16'h00a6,16'h005d,-16'h00ff,-16'h006d,-16'h017b,16'h00d7,-16'h006b,-16'h022f,16'h00c0,16'h00ea,-16'h0057,16'h0277,-16'h0064,-16'h006c,-16'h00a3,16'h0069,16'h0125,-16'h0074,-16'h0079,-16'h003b,16'h015d,-16'h00e8,-16'h00f2,16'h000c,-16'h0079,-16'h0115,16'h0021,16'h0062,-16'h000e,16'h0089,-16'h0236,16'h000d,16'h0033,16'h0274,-16'h0129,16'h0100,-16'h019c,-16'h006f,16'h002d,-16'h0029,16'h00ef,-16'h0156,16'h004b,-16'h0051,-16'h0085,-16'h0019,16'h013c,-16'h0095,-16'h0039,16'h0008,16'h0054,-16'h00e9,16'h0049,16'h0129,16'h017d,16'h000c,16'h00a8,16'h00d8,-16'h0085,-16'h00b5,-16'h0086,16'h002e,-16'h0039,16'h019c,-16'h00c5,16'h00c4,-16'h00dc,-16'h0074,-16'h0150,16'h00f4,-16'h0059,-16'h0168,16'h00ef,16'h00a0,-16'h0085,16'h01d5,-16'h00a6,-16'h00ad,-16'h008e,16'h0040,16'h020c,16'h0001,-16'h0033,16'h0074,-16'h0043,-16'h0084,-16'h0052,-16'h0013,-16'h00a9,-16'h0062,16'h002d,16'h00c5,-16'h0003,16'h0021,-16'h018a,16'h0012,16'h00cd,16'h0242,-16'h024a,16'h008d,-16'h015a,16'h00de,16'h0001,16'h0071,16'h009c,-16'h0150,-16'h004a,-16'h00da,16'h0004,16'h0016,16'h0179,-16'h00cb,16'h0022,-16'h00b1,16'h0070,-16'h00ac,16'h00c3,16'h00dd,16'h0183,-16'h000a,16'h00a4,16'h00bc,-16'h0075,-16'h00db,-16'h00a7,-16'h0026,-16'h0060,16'h0260,-16'h010e,16'h0102,-16'h0056,-16'h005f,-16'h00c3,16'h00da,16'h002c,-16'h0101,16'h0110,16'h007c,-16'h009c,16'h0184,-16'h003d,-16'h0067,-16'h00c9,-16'h0068,16'h0179,-16'h013c,-16'h0001,-16'h005a,-16'h018b,16'h00a2,-16'h005b,-16'h0030,-16'h0131,-16'h00a3,16'h0094,16'h0163,-16'h0027,16'h00dc,-16'h00b6,16'h001a,16'h00ef,16'h01ea,-16'h020c,16'h003b,-16'h00b3,16'h0094,16'h0035,16'h0020,16'h011e,-16'h0074,16'h0012,-16'h006b,16'h0023,16'h0091,16'h00ec,-16'h0072,16'h00c0,-16'h0091,16'h002f,-16'h00ee,16'h0161,16'h0100,16'h0158,16'h0030,16'h001f,16'h00e5,16'h0030,-16'h0118,-16'h0070,-16'h005c,-16'h00fa,16'h01fa,-16'h015f,16'h0173,16'h0005,16'h001a,-16'h0022,16'h0115,16'h00ba,-16'h00e2,16'h0151,16'h003b,-16'h001e,16'h0234,-16'h003e,-16'h0040,-16'h00a7,16'h0051,16'h01a2,-16'h017c,-16'h005a,-16'h00a4,-16'h027c,16'h00fd,16'h0059,16'h001b,-16'h0149,-16'h00ae,16'h0045,16'h00e2,-16'h0006,16'h0000,-16'h005d,-16'h0045,16'h0100,16'h0209,-16'h0175,16'h0032,16'h0049,16'h0111,16'h00d8,16'h0066,16'h00ec,16'h0091,-16'h0013,-16'h005b,16'h0100,-16'h0037,16'h00dd,-16'h009a,16'h007c,-16'h0009,-16'h00b3,-16'h0003,16'h01fe,16'h00cc,16'h01af,-16'h0003,16'h007b,16'h018f,16'h002d,-16'h004e,-16'h0087,-16'h00dc,-16'h0177,16'h0157,-16'h0110,16'h017c,-16'h0158,-16'h0022,-16'h002d,16'h0112,16'h012b,-16'h003d,16'h0116,16'h0026,16'h0093,16'h0218,-16'h0020,-16'h004b,16'h00d4,-16'h001b,16'h0197,-16'h014d,-16'h0029,-16'h008b,-16'h021e,16'h023e,16'h00d4,16'h002e,-16'h017b,-16'h0043,-16'h003d,16'h001e,-16'h00e6,16'h0004,-16'h0048,-16'h00d3,16'h0094,16'h0207,-16'h00d4,16'h006c,16'h00eb,16'h0140,16'h0161,16'h0044,16'h0078,16'h016b,16'h003f,-16'h00af,16'h00aa,-16'h0031,16'h00ed,-16'h0055,16'h0009,16'h0000,-16'h015b,16'h0078,16'h024a,16'h00c2,16'h0152,16'h007a,16'h009a,16'h0098,16'h0039,-16'h0074,-16'h00d9,-16'h008e,-16'h0132,-16'h017a,-16'h005f,16'h0177,-16'h0199,-16'h0012,-16'h0085,16'h00aa,16'h0100,16'h0063,16'h011c,16'h0022,16'h00d2,16'h01ed,16'h0053,-16'h0060,16'h00d1,-16'h0090,16'h00b4,-16'h0159,-16'h00b5,-16'h0089,-16'h0108,16'h016e,16'h010b,16'h0044,-16'h01c7,-16'h003b,-16'h00ff,-16'h00ff,-16'h00f6,-16'h00e9,16'h000e,-16'h00f6,16'h006c,16'h01ea,-16'h00f5,16'h00c3,16'h0085,16'h01ff,16'h00d4,-16'h0036,16'h004c,16'h00fc,16'h00cd,-16'h00c8,16'h00de,-16'h007d,16'h0082,-16'h0075,16'h00b7,-16'h0009,-16'h011d,16'h000a,16'h017d,16'h00d1,16'h01a9,16'h0096,16'h00b9,-16'h0049,16'h0063,-16'h0042,-16'h0052,-16'h00aa,-16'h01be,-16'h02b6,16'h0001,16'h010a,-16'h0056,16'h0039,-16'h00d6,16'h0070,16'h0113,16'h00a2,16'h0100,-16'h0046,16'h010b,16'h0240,16'h0084,-16'h0064,16'h016b,-16'h002d,-16'h0080,-16'h00a9,-16'h00b0,-16'h00ae,-16'h0063,-16'h012d,16'h01da,16'h00aa,-16'h01bf,-16'h0065,-16'h007b,-16'h0056,-16'h0089,-16'h00a1,-16'h00a1,-16'h011a,16'h0034,16'h01ec,-16'h00ac,16'h00c3,16'h00d2,16'h021a,16'h0041,-16'h007c,-16'h0062,16'h00de,16'h011f,-16'h0112,16'h00b5,-16'h0090,16'h00a0,-16'h003e,16'h0017,16'h001e,-16'h0198,16'h00b3,16'h0190,16'h008e,16'h00e1,16'h00b1,16'h0091,-16'h008f,16'h0099,-16'h008f,16'h0031,-16'h0028,-16'h0160,-16'h0168,-16'h0011,16'h00bd,16'h002f,16'h0025,-16'h00d0,16'h00d3,16'h0157,16'h00cf,16'h0148,-16'h0020,16'h002d,16'h01cb,16'h00ce,-16'h0035,-16'h004f,16'h0040,-16'h00bd,16'h0049,-16'h006f,-16'h008a,16'h009a,-16'h033e,16'h0208,16'h00af,-16'h01f4,-16'h004e,16'h001a,-16'h003a,-16'h015d,-16'h00c3,-16'h011e,-16'h00f6,-16'h002d,16'h01e6,16'h00a8,16'h0094,16'h00de,16'h0202,16'h0069,16'h000f,-16'h00f4,16'h005e,16'h0158,-16'h005c,16'h0010,-16'h005f,16'h0037,-16'h0054,-16'h0014,16'h00ce,-16'h01c3,16'h0073,16'h012d,16'h011c,16'h0056,16'h00e6,16'h0139,-16'h00c0,16'h008e,-16'h002b,16'h00e3,-16'h003a,-16'h01ae,-16'h002d,16'h00dd,16'h0129,16'h00b1,-16'h0011,-16'h00eb,16'h001a,16'h005e,16'h0125,16'h006b,16'h009b,-16'h0011,16'h0125,16'h00c1,-16'h0099,-16'h0185,16'h00dc,-16'h0166,16'h00c6,-16'h003d,-16'h0028,16'h0023,-16'h01c1,16'h01cc,16'h016f,-16'h01f3,-16'h00f7,16'h0097,-16'h0050,-16'h018c,16'h0037,-16'h002e,-16'h004b,-16'h006a,16'h0203,16'h00df,16'h00c2,16'h0109,16'h016c,16'h004d,16'h0022,-16'h014c,-16'h00c0,16'h01cb,-16'h003c,16'h0039,-16'h0051,16'h009d,-16'h0097,-16'h010d,16'h005a,-16'h0225,16'h0092,16'h015c,16'h0063,16'h00cb,16'h0163,16'h015b,-16'h0113,16'h00e1,-16'h0001,16'h01a1,16'h003d,-16'h01a0,-16'h0058,16'h013f,16'h0115,16'h007e,-16'h000d,-16'h00da,16'h00e9,-16'h0093,16'h00f1,16'h002e,16'h00ed,-16'h0020,16'h013d,16'h011a,-16'h0067,-16'h0264,16'h00a9,-16'h014b,16'h0151,-16'h0082,-16'h0030,-16'h00a4,16'h011c,16'h0216,16'h0139,-16'h01cd,-16'h00bc,16'h00b2,-16'h00ed,-16'h0170,16'h0092,16'h0049,-16'h002f,-16'h0085,16'h01ac,16'h013b,16'h00ed,16'h0074,16'h0153,16'h002d,16'h008a,-16'h0148,-16'h015f,16'h01a0,-16'h005a,16'h0017,16'h0009,16'h00ad,-16'h00d6,-16'h0114,16'h00a6,-16'h033c,16'h007d,16'h01aa,16'h0079,16'h0044,16'h005c,16'h0174,-16'h00fe,16'h00f5,-16'h0091,16'h01db,16'h0014,-16'h0167,16'h0012,16'h0156,16'h013c,16'h009f,16'h006a,-16'h00bf,16'h0061,-16'h03a1,16'h00d6,-16'h002e,16'h00ca,16'h0014,16'h00ef,16'h00c3,-16'h00c8,-16'h021d,16'h005b,-16'h01da,16'h00b6,-16'h00e2,16'h0045,-16'h004f,16'h0194,16'h0235,-16'h008e,-16'h0251,-16'h00d0,16'h006f,-16'h0067,-16'h00a2,16'h0087,-16'h000a,-16'h0010,-16'h00e8,16'h00f7,16'h0124,16'h0079,16'h009b,16'h01a1,16'h005d,16'h006d,-16'h0040,-16'h0203,16'h01cb,16'h0027,16'h0008,-16'h0078,16'h0075,-16'h00ed,-16'h00f6,16'h00b1,-16'h0420,16'h0094,16'h018d,16'h00da,-16'h004a,16'h004b,16'h0177,-16'h00cf,16'h0149,-16'h001f,16'h0171,16'h0014,-16'h0090,16'h0036,16'h006a,16'h00d7,-16'h000b,16'h0029,-16'h00b1,16'h0045,-16'h0728,16'h003b,-16'h0064,16'h0006,16'h0079,16'h00d3,16'h00d9,-16'h0040,-16'h0144,16'h0036,-16'h0213,16'h0042,-16'h0092,16'h0132,-16'h004f,16'h0151,16'h0226,-16'h02cf,-16'h024e,-16'h0131,-16'h000f,-16'h0096,-16'h0092,16'h004f,-16'h0035,16'h0063,-16'h00b2,16'h015e,16'h00e2,16'h003d,16'h003d,16'h0159,16'h0002,16'h00a5,-16'h0034,-16'h018e,16'h0285,16'h0050,16'h009b,-16'h0025,16'h005e,-16'h0124,-16'h008c,16'h002a,-16'h0517,16'h0060,16'h00f4,16'h008d,-16'h0047,16'h0050,16'h0131,-16'h0002,16'h0095,-16'h0030,16'h00a8,16'h006c,-16'h007f,-16'h0021,-16'h012c,16'h00ed,-16'h006c,16'h0034,-16'h00d0,16'h00c8,-16'h0655,-16'h000a,-16'h007e,-16'h0083,16'h0004,16'h019c,16'h0029,-16'h0082,16'h0136,16'h002a,-16'h0292,-16'h008c,-16'h0033,16'h0182,-16'h0040,16'h0155,16'h0291,-16'h0298,-16'h0233,-16'h01ed,16'h0026,16'h0089,-16'h0036,-16'h003b,-16'h00af,16'h00da,-16'h0126,16'h01ab,16'h00a2,16'h001a,16'h0070,16'h0129,16'h004c,16'h00d7,16'h0067,-16'h00a0,16'h029d,16'h000a,16'h00eb,16'h0054,16'h006a,-16'h00c0,16'h001a,16'h0060,-16'h062f,16'h0024,16'h007b,16'h00f9,-16'h000c,16'h0048,16'h01b7,-16'h003e,16'h0095,16'h002a,16'h004c,16'h0054,16'h006f,-16'h0020,-16'h02f4,16'h00d3,-16'h01f0,-16'h008e,-16'h008e,16'h0031,-16'h040e,16'h0001,-16'h0054,-16'h004e,16'h004d,16'h0246,16'h006a,-16'h0030,16'h01cd,-16'h002a,-16'h01e5,-16'h0192,16'h0089,16'h01f0,16'h0023,-16'h004c,16'h0231,-16'h01d7,-16'h01ba,-16'h018a,16'h003f,16'h0072,-16'h006f,-16'h010c,-16'h00aa,16'h0168,-16'h0186,16'h00e2,-16'h0006,16'h0022,-16'h0024,16'h012f,16'h00c6,16'h00ba,16'h00cb,16'h0017,16'h01f4,16'h0018,16'h00f6,16'h005a,16'h00e0,-16'h0144,16'h0140,16'h00a2,-16'h05e6,16'h00c9,16'h008b,16'h00b9,-16'h0033,16'h007a,16'h015a,-16'h00b9,16'h00c8,16'h0040,-16'h002c,16'h0089,16'h002e,16'h000d,-16'h0628,16'h0070,-16'h029b,-16'h007b,-16'h00b3,-16'h0033,-16'h025c,-16'h00e7,-16'h0038,-16'h0004,16'h006e,16'h017b,16'h003b,-16'h009b,16'h01b4,-16'h00f9,-16'h0095,-16'h0138,16'h0057,16'h0184,-16'h0006,-16'h01b5,16'h02a2,16'h002e,-16'h011f,-16'h0155,16'h00cc,16'h00f0,16'h0069,-16'h02dc,-16'h00d2,16'h0095,-16'h0147,16'h00db,-16'h0020,-16'h0007,-16'h00e9,16'h00f8,16'h005c,-16'h00ac,16'h00aa,-16'h001c,16'h013a,-16'h002e,16'h0183,16'h0074,16'h0029,-16'h011b,16'h014e,16'h00ea,-16'h04ef,16'h0031,16'h0033,16'h0077,-16'h007b,16'h012c,16'h01d6,-16'h0207,16'h00e3,16'h010a,-16'h0081,16'h0045,16'h0042,16'h0053,-16'h056e,16'h000c,-16'h0184,-16'h00cf,-16'h0071,-16'h001c,-16'h019a,-16'h003d,16'h0019,-16'h003a,16'h003a,16'h00b2,16'h0077,-16'h00a6,16'h005e,-16'h009e,-16'h005f,-16'h016f,16'h0012,16'h0105,16'h0098,-16'h024b,16'h0280,16'h01af,-16'h006e,-16'h0150,16'h00a5,16'h0133,16'h00d0,-16'h0475,-16'h012b,16'h0060,-16'h00c7,16'h00d5,16'h0022,-16'h0089,-16'h0167,16'h005a,16'h0004,-16'h00d4,16'h0162,16'h002c,16'h01be,-16'h00a7,16'h0187,16'h00c0,-16'h0081,-16'h010e,16'h00a4,16'h0108,-16'h04af,-16'h007e,16'h0008,16'h00c8,-16'h007b,16'h0107,16'h018c,-16'h0374,16'h0090,16'h0124,-16'h00bf,16'h0036,-16'h0027,16'h0075,-16'h036f,-16'h0029,-16'h00d0,-16'h00fa,-16'h0066,-16'h000f,-16'h00eb,-16'h0068,-16'h000c,-16'h0053,-16'h000d,16'h00ba,-16'h004f,-16'h00c3,-16'h00c7,-16'h00ab,16'h001b,-16'h00d9,-16'h015f,-16'h0088,-16'h0006,-16'h005e,16'h02f3,16'h02fc,-16'h0073,-16'h01d4,16'h00db,16'h0138,16'h0059,-16'h03fc,-16'h01ec,16'h0017,-16'h005b,16'h0162,16'h002a,16'h006c,-16'h00b5,-16'h000a,-16'h0028,-16'h0106,16'h01b5,16'h002e,16'h00c9,-16'h00d9,16'h0000,16'h0040,-16'h006a,-16'h0065,16'h00d3,16'h0060,-16'h041e,-16'h0148,-16'h002e,16'h003d,-16'h00b8,16'h00b6,16'h01d0,-16'h02e8,16'h00be,16'h014a,-16'h014c,16'h0130,-16'h005a,-16'h000c,-16'h00ca,16'h0009,16'h00b4,-16'h00c6,-16'h0045,16'h0058,-16'h009e,16'h0033,-16'h0008,-16'h001d,16'h0002,16'h00f5,-16'h0063,-16'h0068,-16'h0151,-16'h01f6,16'h0044,-16'h0137,-16'h02ef,-16'h00dd,-16'h004a,16'h006e,16'h027d,16'h02af,16'h0015,-16'h014c,16'h00fb,16'h0196,16'h0106,-16'h02da,-16'h02d3,-16'h00d6,16'h0012,16'h011f,16'h00d0,16'h00b2,-16'h0073,16'h0063,-16'h0062,-16'h013f,16'h01e4,-16'h0040,16'h012f,-16'h007c,-16'h025a,-16'h0085,-16'h004e,-16'h004f,16'h008e,16'h00e4,-16'h0324,-16'h0116,-16'h0062,16'h001b,-16'h0096,16'h00cf,16'h0165,-16'h021b,16'h0175,16'h0190,-16'h0203,16'h00b7,16'h0001,-16'h0037,16'h018f,-16'h00c0,16'h01f9,-16'h006c,-16'h00dd,16'h0090,-16'h0048,-16'h0056,-16'h004b,16'h009b,16'h0067,16'h00a3,-16'h0042,-16'h0023,-16'h0114,-16'h01e4,16'h0021,-16'h0007,-16'h0407,-16'h00a0,-16'h00e4,16'h0076,16'h02d2,16'h01f2,-16'h0025,-16'h0155,16'h00e2,16'h0232,16'h00a1,-16'h029b,-16'h0235,-16'h0104,16'h00de,16'h015c,16'h00e6,16'h0071,-16'h010e,-16'h0090,-16'h001b,-16'h0113,16'h017d,-16'h00ac,16'h0106,-16'h006c,-16'h0215,16'h0073,-16'h009f,-16'h0012,16'h00a2,16'h003c,-16'h0247,-16'h015f,-16'h0172,-16'h00c2,-16'h0127,16'h0126,16'h012d,-16'h0128,16'h013a,16'h00e2,-16'h0321,16'h015f,16'h00bd,16'h0016,16'h02a1,-16'h007e,16'h01d1,16'h0041,-16'h0100,16'h0175,-16'h0095,-16'h0040,-16'h00bb,16'h0049,-16'h00ce,16'h00d8,16'h004a,-16'h00e7,-16'h004b,-16'h00c6,16'h00bc,-16'h0006,-16'h0307,16'h0029,-16'h001a,16'h009b,16'h039a,16'h00f0,16'h0041,-16'h00b9,16'h0135,16'h0335,16'h009e,-16'h0179,-16'h01d8,-16'h00b5,16'h0156,16'h0145,16'h003d,16'h00da,-16'h0186,-16'h00d0,-16'h00b0,-16'h0064,16'h0176,-16'h006f,16'h00f6,-16'h00f0,-16'h020e,16'h0143,-16'h010d,-16'h008b,-16'h004a,16'h0161,-16'h01c0,-16'h0068,-16'h0091,16'h001f,-16'h017b,-16'h001a,16'h016b,-16'h00f4,16'h000e,-16'h002a,16'h0054,16'h013c,-16'h005f,16'h00c7,16'h00db,16'h0114,-16'h00a0,-16'h00c4,16'h0076,-16'h0091,16'h0045,16'h0035,16'h0102,16'h00b9,-16'h0010,16'h01da,16'h0023,-16'h0076,-16'h005c,16'h0047,16'h0010,-16'h005e,-16'h009a,-16'h00fe,16'h00a0,-16'h0075,-16'h009c,16'h00bc,16'h0040,16'h00f7,-16'h01aa,16'h0061,16'h001b,16'h0188,-16'h0115,-16'h004f,16'h0064,-16'h000b,16'h0078,16'h007f,-16'h0042,-16'h0111,16'h001c,-16'h0090,16'h00b1,16'h0150,16'h0117,16'h0076,-16'h004f,-16'h0096,16'h0082,16'h00bd,16'h008f,16'h017e,-16'h01b5,-16'h00ab,-16'h0082,16'h00ff,-16'h014b,16'h0035,16'h0109,-16'h015d,16'h0009,16'h00bd,-16'h007b,16'h0186,-16'h0072,16'h0057,-16'h003d,16'h00f0,16'h0019,-16'h00a1,16'h0035,-16'h0062,16'h000e,-16'h00a3,-16'h0070,-16'h0049,-16'h0087,16'h01b3,-16'h004c,-16'h0024,-16'h0070,16'h0056,-16'h0094,-16'h00be,-16'h00e5,-16'h0039,16'h0024,-16'h0022,-16'h00cf,16'h003b,16'h0060,16'h011d,-16'h0198,-16'h0016,16'h00ef,16'h00df,-16'h0155,-16'h0021,16'h0030,16'h0071,16'h00a8,16'h010c,-16'h0160,-16'h0083,16'h0014,16'h0035,16'h00ed,16'h00fc,16'h00b4,16'h0080,-16'h000f,-16'h008f,16'h003b,16'h0025,16'h0012,16'h00da,-16'h00f9,-16'h0118,-16'h010f,16'h00ef,-16'h015e,16'h005b,16'h00da,-16'h0180,16'h0054,16'h00c8,-16'h00c4,16'h008a,16'h0015,16'h01aa,-16'h0035,16'h0139,-16'h0047,-16'h00a6,16'h00a0,16'h009f,16'h0079,-16'h0290,-16'h00c3,-16'h0034,16'h0072,16'h0122,-16'h0065,16'h000e,-16'h0050,16'h0011,-16'h0045,-16'h00cb,-16'h00c1,16'h0057,-16'h004b,16'h001c,-16'h00b5,16'h002b,16'h0027,16'h012d,-16'h018f,-16'h0004,16'h013a,16'h00e2,-16'h0168,-16'h0064,16'h0072,16'h00b1,16'h00c2,16'h00cb,-16'h0125,-16'h012f,-16'h0003,16'h009e,16'h0097,16'h0143,16'h00e3,16'h00c1,16'h005a,-16'h007f,-16'h00a9,16'h0011,-16'h008b,16'h007c,-16'h00bd,-16'h0045,-16'h00cc,16'h00b4,-16'h00c1,16'h0057,16'h00cd,-16'h00df,16'h002d,16'h0068,-16'h00f2,16'h0089,-16'h002e,16'h015d,-16'h0055,16'h00cc,-16'h00b5,-16'h0041,16'h0073,16'h0119,16'h00a0,-16'h02f7,-16'h00e0,-16'h007b,16'h004e,16'h017c,-16'h0040,-16'h006f,16'h0013,16'h007b,16'h0036,16'h000b,-16'h00f3,16'h0060,-16'h0049,-16'h0033,-16'h0086,-16'h0036,-16'h000a,16'h012e,-16'h0120,16'h003b,16'h0084,16'h00ee,-16'h01fa,-16'h0080,16'h0048,16'h00fa,16'h012a,16'h00c4,-16'h0185,-16'h00b0,-16'h002e,16'h0029,16'h00af,16'h017a,16'h013d,16'h00d2,16'h008c,-16'h0048,-16'h002f,-16'h002e,-16'h0112,16'h00c3,-16'h0063,-16'h0076,-16'h00a6,16'h0155,-16'h0085,-16'h004c,16'h00ac,-16'h003a,16'h0007,-16'h0050,-16'h0086,16'h00f7,-16'h0045,16'h0056,-16'h009d,16'h0132,-16'h000d,-16'h003c,16'h003d,16'h0063,16'h0040,-16'h01bc,-16'h02bf,-16'h003e,16'h009a,16'h0224,16'h003a,-16'h0097,16'h0050,16'h0090,16'h009b,16'h0038,-16'h0115,16'h000d,-16'h00a6,-16'h0099,-16'h0095,16'h0054,-16'h0006,16'h0146,-16'h007b,-16'h0073,16'h0086,16'h006b,-16'h0264,-16'h0056,16'h005a,16'h01dd,16'h0145,16'h00f4,-16'h01b0,-16'h010f,16'h0006,-16'h002e,16'h0116,16'h013d,16'h0108,16'h00d6,16'h0012,-16'h00be,-16'h0128,16'h000c,-16'h01ba,16'h00c4,16'h00b0,16'h0003,-16'h00d4,16'h0133,-16'h00ea,-16'h0012,16'h00f4,16'h014e,-16'h0032,-16'h0042,16'h0013,16'h00ed,-16'h0059,-16'h012b,-16'h0023,16'h015e,-16'h0071,-16'h0079,-16'h0025,16'h00b9,16'h002b,-16'h0147,-16'h0419,16'h004d,16'h004e,16'h0285,16'h0058,-16'h0017,-16'h0010,16'h005a,16'h00a6,-16'h0046,-16'h00d4,-16'h001d,-16'h0048,-16'h006d,-16'h0030,16'h0070,-16'h0077,16'h0043,16'h001a,-16'h000c,-16'h0079,16'h0114,-16'h030a,16'h000f,16'h0007,16'h01f5,16'h019c,16'h0135,-16'h01e3,-16'h017a,16'h0038,-16'h0009,16'h00c4,16'h00a3,16'h0061,16'h0062,-16'h006f,-16'h0024,-16'h008a,-16'h0090,-16'h0125,16'h0085,16'h00f9,-16'h00b6,-16'h00e4,16'h0164,-16'h0024,16'h002c,16'h00c8,16'h0185,-16'h0037,-16'h0083,16'h005f,16'h0085,-16'h0054,-16'h0382,-16'h004e,16'h00e5,-16'h0024,-16'h00a6,16'h0001,-16'h0026,16'h0023,-16'h0112,-16'h020b,16'h0009,16'h0033,16'h0273,16'h0047,-16'h00a0,-16'h00a0,16'h0094,16'h00e4,-16'h001c,-16'h0061,-16'h00be,16'h00ed,-16'h008f,-16'h00ed,-16'h0009,-16'h0078,-16'h003a,-16'h0029,16'h0007,-16'h0053,16'h00e6,-16'h02e2,16'h002c,16'h0092,16'h026f,16'h011c,16'h0195,-16'h0132,-16'h0218,16'h0159,-16'h004a,16'h00e0,-16'h0036,16'h0055,16'h0018,-16'h00d1,-16'h0053,-16'h000c,-16'h0090,-16'h0051,16'h0053,16'h00c0,-16'h01b2,-16'h00a8,16'h0128,16'h002e,-16'h0044,16'h00f7,16'h01c0,-16'h0040,-16'h00b0,16'h003c,-16'h0010,16'h0091,-16'h0236,-16'h006e,16'h012f,16'h0001,-16'h006e,16'h0046,16'h002a,-16'h0084,-16'h01fa,16'h007f,16'h00ce,16'h001a,16'h0265,-16'h0015,-16'h008c,-16'h00c1,16'h00df,16'h0173,-16'h006a,-16'h0047,-16'h0036,16'h01bd,-16'h0137,-16'h00c7,16'h0023,-16'h00d9,-16'h0033,-16'h003c,16'h00c1,-16'h006f,16'h00d1,-16'h0210,16'h004d,16'h00dc,16'h02a4,-16'h001f,16'h0144,-16'h01a9,-16'h02c1,16'h00df,-16'h004e,16'h00eb,-16'h0171,16'h004d,-16'h001f,-16'h003f,-16'h0012,16'h00a5,-16'h0099,-16'h0012,-16'h005b,-16'h0002,-16'h01a2,-16'h0007,16'h015a,16'h00f4,-16'h008d,16'h0123,16'h0148,-16'h0057,-16'h00fa,16'h0098,-16'h0008,16'h0079,16'h0037,-16'h0091,16'h00ce,-16'h002b,16'h000a,-16'h008e,16'h0063,-16'h0050,-16'h01ab,16'h00d2,16'h010a,-16'h0008,16'h0232,-16'h0045,-16'h0020,-16'h00e7,16'h00bb,16'h017b,-16'h0089,-16'h0012,16'h008f,16'h0140,-16'h00f7,-16'h009f,16'h0017,-16'h00a5,-16'h004c,-16'h00a9,16'h0073,-16'h0087,16'h00a2,-16'h018d,16'h0044,16'h00da,16'h02b0,-16'h01b6,16'h00e3,-16'h019d,-16'h0344,16'h0061,16'h003e,16'h0099,-16'h01d7,-16'h0050,-16'h00a3,-16'h001b,-16'h0068,16'h00a9,-16'h00c1,16'h006e,-16'h006b,16'h0031,-16'h0132,16'h00dd,16'h0098,16'h011a,-16'h003d,16'h006d,16'h0158,-16'h0049,-16'h00fe,16'h0009,-16'h0066,16'h0014,16'h0267,-16'h003e,16'h00d1,-16'h0036,-16'h0053,-16'h0065,16'h0073,-16'h0052,-16'h0107,16'h014a,16'h0043,-16'h0107,16'h01f3,-16'h009b,-16'h0089,-16'h006c,16'h00b1,16'h01b9,-16'h013b,-16'h0065,16'h0067,-16'h006e,-16'h0093,-16'h00b3,-16'h0036,-16'h0109,16'h0025,-16'h005f,16'h00a8,16'h0002,16'h003f,-16'h0039,16'h0020,16'h00d3,16'h021f,-16'h0200,16'h00ba,-16'h00e3,-16'h0382,16'h0019,16'h00e2,16'h005e,-16'h00c6,-16'h009e,-16'h00fe,16'h0026,16'h000b,16'h012d,-16'h00b7,16'h00c1,-16'h00c7,16'h0008,-16'h012f,16'h0123,16'h0177,16'h014c,-16'h0017,16'h0055,16'h0009,-16'h0006,-16'h017a,-16'h0081,-16'h00bc,16'h0073,16'h0233,-16'h00b1,16'h0135,16'h0086,-16'h00a8,-16'h0057,16'h002d,-16'h00a6,-16'h0069,16'h0184,16'h0030,-16'h00c0,16'h0138,-16'h0085,-16'h0080,-16'h0055,16'h005a,16'h01a4,-16'h01e3,-16'h0059,-16'h0054,-16'h0243,16'h0062,-16'h00f9,16'h0090,-16'h0095,-16'h0046,16'h0036,16'h0151,16'h001b,16'h0059,-16'h0027,16'h0011,16'h00dd,16'h028c,-16'h019f,16'h00b9,16'h0031,-16'h032e,16'h00d8,16'h0078,16'h002a,16'h005c,-16'h0041,-16'h00c3,16'h0089,-16'h0012,16'h0161,-16'h00fe,16'h0120,-16'h0094,-16'h003c,-16'h00fb,16'h014f,16'h0109,16'h0190,-16'h003b,16'h0015,16'h00b4,16'h0009,-16'h00d1,-16'h005f,-16'h0051,16'h0002,16'h0160,-16'h0098,16'h00e4,-16'h002b,-16'h0042,-16'h0002,16'h004d,16'h0027,16'h001a,16'h014e,16'h0041,16'h0042,16'h01f1,-16'h008a,-16'h003f,-16'h0084,16'h0021,16'h023c,-16'h01c3,-16'h007b,-16'h0043,-16'h0306,16'h0146,-16'h00c4,16'h0003,-16'h011e,-16'h00d2,16'h004e,16'h0194,16'h0015,16'h001a,16'h003e,-16'h0055,16'h0140,16'h0223,-16'h00dc,16'h00ac,16'h00a5,-16'h02f7,16'h017e,16'h0037,16'h0014,16'h00f3,-16'h0015,-16'h0076,16'h009c,-16'h0014,16'h0185,-16'h00c4,16'h0130,-16'h0002,-16'h0119,-16'h00bd,16'h0151,16'h012f,16'h0177,16'h0095,16'h00a7,16'h00d3,16'h0085,-16'h000f,-16'h0123,-16'h00b2,-16'h0078,16'h0069,-16'h00d2,16'h0179,-16'h00b4,-16'h0090,16'h0036,16'h001a,16'h00c1,16'h006b,16'h0127,-16'h0007,16'h0105,16'h023e,-16'h0079,-16'h00fc,16'h006c,-16'h0085,16'h018e,-16'h0182,-16'h0069,-16'h0003,-16'h016d,16'h0252,-16'h00c4,-16'h005e,-16'h0153,16'h000f,-16'h00b0,16'h009e,-16'h0078,-16'h0075,16'h0075,-16'h00bb,16'h00ee,16'h01c8,-16'h00e1,16'h008c,16'h00b9,-16'h0244,16'h0101,16'h003e,-16'h0003,16'h01ce,16'h0029,-16'h00b4,16'h00e2,-16'h0020,16'h00f3,-16'h00d5,16'h0092,-16'h0039,-16'h00e7,16'h002b,16'h01a3,16'h016c,16'h01a5,16'h0019,16'h00d7,16'h0052,16'h006d,16'h006a,-16'h006e,-16'h0108,-16'h00d1,-16'h01ca,-16'h00d3,16'h0114,-16'h00c5,-16'h0031,-16'h00b4,16'h00a8,16'h0168,16'h00dd,16'h00a0,16'h0046,16'h01a4,16'h01fc,16'h0061,-16'h00fd,16'h00ee,-16'h00e2,16'h00c1,-16'h00a1,-16'h009d,-16'h004d,-16'h006f,16'h011a,-16'h000e,-16'h003c,-16'h0103,-16'h005c,-16'h0091,-16'h0058,16'h0012,-16'h0099,16'h0010,-16'h0143,16'h0087,16'h016d,-16'h0112,16'h008e,16'h00d6,-16'h01ea,16'h015a,-16'h0001,-16'h002c,16'h01ab,16'h0011,-16'h00b7,16'h00c8,-16'h003f,16'h00fc,-16'h00a2,16'h0007,-16'h0025,-16'h0074,-16'h004f,16'h0163,16'h0158,16'h0114,16'h0024,16'h00fa,-16'h00a2,16'h00db,16'h000c,-16'h0016,-16'h0130,-16'h00f9,-16'h0272,-16'h00ac,16'h00a6,-16'h0002,16'h0046,-16'h00dd,16'h00d4,16'h01da,-16'h0010,16'h00c3,16'h0001,16'h01cb,16'h0225,16'h0033,-16'h00a7,16'h00e7,-16'h0052,-16'h00b4,16'h0035,-16'h00bb,-16'h00a2,16'h0003,-16'h0289,16'h0008,16'h0040,-16'h00ed,-16'h00f7,-16'h0047,-16'h00a0,-16'h0097,-16'h005e,16'h0038,-16'h012b,16'h012b,16'h0174,-16'h00a7,16'h0061,16'h011b,-16'h01d6,16'h010a,16'h0048,-16'h004a,16'h00cc,16'h0140,-16'h005b,16'h0046,16'h0045,16'h0100,-16'h00d7,16'h0020,16'h0020,-16'h0131,16'h0008,16'h0196,16'h0155,16'h0195,16'h0089,16'h009f,-16'h00a2,16'h00fc,16'h002f,16'h0022,-16'h007c,-16'h0146,-16'h0088,-16'h0025,16'h00c9,16'h007d,16'h0059,-16'h0115,16'h0120,16'h01a0,16'h00d0,16'h000d,-16'h0027,16'h00f8,16'h01fe,16'h008c,-16'h00c2,16'h004b,16'h0048,-16'h00f1,16'h00e6,-16'h00d9,-16'h0102,16'h0094,-16'h0450,16'h00d1,16'h00b1,-16'h0148,-16'h015f,16'h0032,-16'h0062,-16'h011a,-16'h0058,16'h000d,-16'h00b2,16'h00ea,16'h01a5,16'h000a,16'h0078,16'h0128,-16'h014d,16'h010e,16'h008a,-16'h00e0,16'h0095,16'h00ef,-16'h008b,-16'h005c,-16'h005c,16'h00a8,-16'h0108,-16'h00db,16'h004d,-16'h007a,16'h0029,16'h00f0,16'h0119,16'h0112,16'h00c1,16'h0128,-16'h010e,16'h00d8,16'h0075,16'h007e,-16'h009b,-16'h018a,16'h0037,16'h004f,16'h00aa,16'h007e,-16'h0004,-16'h012f,16'h00b6,16'h0113,16'h0086,-16'h007e,16'h006c,-16'h0042,16'h0118,16'h0133,-16'h0090,-16'h0137,16'h0105,-16'h0114,16'h0103,-16'h0076,-16'h0134,16'h000d,-16'h016d,16'h010a,16'h0111,-16'h018d,-16'h0075,16'h00a7,-16'h0094,-16'h0137,-16'h0062,-16'h0042,-16'h0065,-16'h0033,16'h01cc,16'h002d,16'h001e,16'h00eb,-16'h0120,16'h00f2,16'h0124,-16'h0158,-16'h00c8,16'h012b,-16'h006b,-16'h0038,-16'h000f,16'h0071,-16'h016a,-16'h0142,16'h0122,-16'h006c,-16'h00a8,16'h010e,16'h00c0,16'h0136,16'h0135,16'h019e,-16'h00c4,16'h0084,16'h0036,16'h0108,-16'h0044,-16'h016a,16'h013b,16'h014b,16'h00af,16'h00c3,16'h001a,-16'h019f,16'h0081,-16'h0033,16'h00f3,-16'h014d,16'h005a,-16'h009d,16'h00d3,16'h0166,-16'h00f4,-16'h0144,16'h0134,-16'h015a,16'h0121,-16'h0194,-16'h011e,-16'h0084,16'h0135,16'h00c3,16'h00f0,-16'h01ba,-16'h0037,16'h0059,-16'h00ee,-16'h0152,16'h001d,-16'h0016,16'h0008,-16'h0093,16'h018f,16'h00c3,16'h0046,16'h00dc,-16'h00a4,16'h0060,16'h013d,-16'h0198,-16'h0166,16'h01cd,-16'h00ab,16'h0007,-16'h005c,16'h0062,-16'h0120,-16'h00d3,16'h0151,-16'h00bc,-16'h0060,16'h01a2,16'h00c2,16'h007e,16'h010b,16'h0138,-16'h0085,16'h00bd,-16'h0003,16'h011e,-16'h005b,-16'h015d,16'h008d,16'h01c3,16'h0046,16'h0111,16'h0043,-16'h015e,16'h0098,-16'h01ed,16'h0091,-16'h0103,16'h0021,-16'h002b,16'h00da,16'h0185,-16'h0119,-16'h01dc,16'h004d,-16'h010c,16'h0097,-16'h00e6,-16'h0057,-16'h0082,16'h0125,16'h00e7,-16'h008e,-16'h0244,16'h0008,16'h00ac,-16'h00ec,-16'h0163,16'h00c9,-16'h0068,16'h0074,-16'h0087,16'h014b,16'h0126,16'h001b,-16'h0004,-16'h00b3,16'h002b,16'h0144,-16'h00dd,-16'h00fd,16'h0156,-16'h005c,16'h0063,-16'h00e5,-16'h0014,-16'h00c7,-16'h00af,16'h0107,-16'h018a,-16'h00c9,16'h0124,16'h0182,16'h0070,16'h00a5,16'h00d8,16'h001d,16'h0192,16'h0006,16'h009c,16'h0043,-16'h011d,16'h00c2,16'h0142,-16'h0007,16'h0055,16'h0066,-16'h00f8,16'h00d0,-16'h05e3,-16'h0002,-16'h0069,-16'h0037,-16'h005c,16'h0160,16'h00b5,-16'h00b3,-16'h0120,16'h005c,-16'h0135,-16'h0038,-16'h008f,16'h0111,16'h000f,16'h0125,16'h019c,-16'h02c9,-16'h019e,16'h001a,16'h000c,-16'h005e,-16'h0138,16'h0000,-16'h00d0,16'h00c0,-16'h00ce,16'h0144,16'h00c9,-16'h004d,-16'h0007,-16'h00a2,16'h0065,16'h00d9,-16'h00a4,-16'h00d1,16'h01eb,-16'h001f,16'h0080,-16'h0004,16'h0016,-16'h011b,-16'h0041,16'h00db,-16'h030a,-16'h0039,16'h015f,16'h016e,16'h008e,16'h0058,16'h011e,16'h0055,16'h0116,16'h001e,16'h00ef,16'h0082,-16'h0074,16'h001c,-16'h00dd,16'h000e,16'h0043,16'h003a,-16'h00d1,16'h006b,-16'h0661,-16'h004c,-16'h00bd,-16'h0061,16'h002e,16'h012a,16'h0041,-16'h00de,16'h00a7,16'h009b,-16'h0076,-16'h00ad,-16'h003b,16'h01a8,16'h0014,16'h013a,16'h0117,-16'h02f1,-16'h0196,-16'h0055,16'h0000,16'h0082,-16'h0130,-16'h0090,-16'h012c,-16'h0002,-16'h0125,16'h00ed,16'h0133,16'h0043,-16'h0073,-16'h0077,16'h009e,16'h0053,16'h0025,-16'h007f,16'h01cd,16'h004b,16'h00b2,-16'h0018,16'h00cf,-16'h00e4,-16'h005c,16'h0037,-16'h0547,-16'h0042,16'h0121,16'h00e4,16'h0010,16'h008f,16'h0170,16'h004f,16'h013d,16'h0096,16'h0042,16'h0065,-16'h0012,-16'h0055,-16'h037b,-16'h000d,-16'h00c8,16'h0006,-16'h0010,-16'h000e,-16'h040a,-16'h0056,-16'h0126,-16'h0032,16'h0058,16'h0193,-16'h0039,-16'h00ea,16'h0151,-16'h0026,-16'h006e,-16'h0110,-16'h0047,16'h0200,16'h0008,-16'h0021,16'h0111,-16'h0185,-16'h018f,-16'h0081,16'h0027,16'h00ef,-16'h0065,16'h007b,-16'h011e,16'h0086,-16'h0127,16'h010b,16'h00a4,16'h007f,-16'h0078,-16'h0012,16'h006c,-16'h0042,16'h00d9,-16'h0007,16'h01af,16'h0012,16'h012f,16'h005e,16'h009f,-16'h015e,16'h0040,16'h005a,-16'h057f,-16'h00bf,16'h011f,16'h00cd,16'h004c,16'h009b,16'h0182,-16'h0031,16'h015c,16'h001d,16'h003c,16'h0001,-16'h0078,-16'h0031,-16'h06a9,-16'h0122,-16'h01c1,-16'h001d,16'h0000,-16'h00b1,-16'h0267,-16'h00b9,-16'h00a4,-16'h0089,16'h002e,16'h01ea,-16'h0122,-16'h00ba,16'h017c,-16'h0015,16'h001e,-16'h00d2,16'h0028,16'h00ee,16'h0001,-16'h01e4,16'h0173,16'h0022,-16'h01bd,-16'h00fc,16'h0008,16'h01bd,-16'h001b,-16'h0118,-16'h0195,16'h0032,-16'h00e5,16'h00f3,16'h005b,16'h0098,-16'h00d2,16'h0029,-16'h0047,-16'h0254,16'h015b,16'h0099,16'h00fd,16'h0000,16'h015b,16'h0019,16'h0020,-16'h012f,16'h00a9,16'h00d9,-16'h0538,-16'h01a5,16'h01f3,16'h00e4,-16'h0072,16'h00fe,16'h01d1,-16'h010a,16'h00ff,16'h00c0,-16'h0037,16'h005d,-16'h0030,-16'h008f,-16'h05d5,-16'h0136,-16'h0180,-16'h0102,16'h0067,-16'h0096,-16'h019a,-16'h0034,-16'h004b,-16'h00c0,16'h004d,16'h0152,-16'h014a,-16'h001d,16'h007b,-16'h00c4,16'h0097,-16'h00af,-16'h0055,16'h0000,16'h0024,-16'h02c0,16'h01f1,16'h01be,-16'h00c4,-16'h00bb,16'h00e2,16'h01bd,16'h002d,-16'h0261,-16'h0221,16'h0011,-16'h0078,16'h013c,16'h0055,16'h00a0,-16'h009d,16'h0082,-16'h00c7,-16'h0248,16'h01af,16'h00e8,16'h00b4,-16'h006e,16'h00b1,16'h0068,16'h001d,-16'h0106,16'h0080,16'h00d0,-16'h0480,-16'h020e,16'h016e,16'h003e,-16'h0071,16'h0123,16'h01e9,-16'h016a,16'h00ea,16'h00c0,-16'h0056,16'h0098,-16'h0073,16'h0001,-16'h03c5,-16'h0090,-16'h0067,-16'h0119,16'h0032,-16'h0024,-16'h00e4,16'h0013,-16'h0089,-16'h009b,16'h0060,16'h0116,-16'h01ca,-16'h0087,-16'h0120,-16'h00db,16'h0078,-16'h009a,-16'h00ea,-16'h0168,-16'h0035,-16'h00e0,16'h0205,16'h033d,-16'h0035,-16'h0139,16'h00ad,16'h01b8,16'h0016,-16'h02b4,-16'h022b,16'h0045,-16'h000f,16'h0112,16'h007f,16'h0099,-16'h0023,16'h0055,-16'h00b6,-16'h0177,16'h0164,16'h0054,16'h00f8,-16'h0106,-16'h011b,16'h0067,-16'h009d,-16'h00a8,16'h0034,16'h00ae,-16'h03c5,-16'h0304,16'h00d2,16'h00b5,-16'h00b9,16'h00a7,16'h016e,-16'h01b0,16'h0144,16'h0154,-16'h00ef,16'h00d0,16'h0047,16'h005c,-16'h0036,-16'h00b6,16'h00e2,-16'h00f6,-16'h0010,16'h00a2,-16'h0075,-16'h0068,-16'h00c5,16'h000d,16'h006c,16'h00e0,-16'h01db,16'h0019,-16'h01ae,-16'h02bf,16'h00f1,-16'h0098,-16'h01fc,-16'h01af,-16'h0071,16'h00c8,16'h0296,16'h021f,-16'h0023,-16'h0173,16'h00df,16'h015e,16'h00d1,-16'h01a9,-16'h023c,-16'h0072,16'h0098,16'h00cc,16'h0074,16'h00c2,-16'h004a,16'h003a,-16'h0063,-16'h00a8,16'h01be,-16'h003f,16'h00df,-16'h0121,-16'h027e,-16'h0020,-16'h004a,-16'h00d3,16'h009d,16'h0111,-16'h0310,-16'h023d,16'h000a,16'h007d,-16'h00d9,16'h00f8,16'h0177,-16'h013d,16'h014e,16'h0157,-16'h01b7,16'h0043,16'h0074,-16'h007d,16'h01c2,-16'h011b,16'h0204,-16'h0106,-16'h009b,16'h00e7,-16'h00bb,-16'h0100,-16'h00ec,16'h00dc,16'h006b,16'h00a1,-16'h00b9,-16'h004b,-16'h009a,-16'h03d7,16'h00e4,-16'h0019,-16'h038c,-16'h016e,-16'h007d,16'h0092,16'h02a3,16'h01a0,-16'h0057,-16'h01e9,16'h019b,16'h0246,16'h011c,-16'h01c6,-16'h023b,-16'h00c4,16'h00c4,16'h00a0,16'h0060,16'h0110,-16'h0127,-16'h000c,16'h003f,-16'h00c5,16'h01bc,16'h000e,16'h0136,-16'h00a5,-16'h021b,16'h000f,-16'h0023,-16'h00af,16'h00c3,16'h00b8,-16'h0237,-16'h0223,-16'h011c,-16'h0055,-16'h014d,16'h00ee,16'h011c,-16'h0134,16'h0181,16'h004c,-16'h02ae,16'h010d,-16'h0005,16'h0079,16'h02c1,-16'h00ec,16'h0263,-16'h0069,-16'h00d2,16'h00eb,-16'h006b,-16'h00e6,-16'h00c1,16'h0124,-16'h0058,16'h00c3,-16'h0029,-16'h00ec,-16'h0027,-16'h026e,16'h011e,-16'h0091,-16'h03c3,-16'h009c,16'h003b,16'h00ed,16'h0344,16'h005c,-16'h00b2,-16'h0134,16'h015f,16'h0325,16'h00a5,-16'h0194,-16'h023f,-16'h006c,16'h0190,16'h00ec,-16'h004a,16'h00a3,-16'h011a,-16'h004c,-16'h0046,-16'h00c3,16'h019d,16'h0025,16'h016a,-16'h0050,-16'h0100,16'h010e,-16'h00f1,-16'h007c,-16'h0012,16'h01b9,-16'h0146,-16'h008c,-16'h00f0,-16'h0043,-16'h0103,-16'h002c,16'h017e,-16'h00af,-16'h0056,16'h002c,16'h000d,16'h026e,-16'h0117,16'h00b7,16'h008c,16'h0148,-16'h0039,-16'h00bf,16'h006e,16'h0043,16'h0110,16'h0056,16'h0069,16'h004f,-16'h00be,16'h018e,16'h0052,-16'h0005,-16'h00a2,-16'h004a,-16'h000c,-16'h0050,-16'h007b,-16'h0085,16'h00d7,-16'h0065,-16'h00cf,16'h0088,-16'h0039,16'h019a,-16'h018e,16'h00b8,16'h006c,16'h013b,-16'h00ef,-16'h0046,16'h008b,-16'h00e6,-16'h0008,16'h0156,16'h0004,-16'h0049,-16'h006c,-16'h00d3,16'h0067,16'h013f,16'h00fa,16'h00e0,-16'h0094,16'h0027,-16'h0008,16'h0103,16'h009b,16'h01c0,-16'h0169,-16'h00b2,-16'h00c7,16'h0027,-16'h01b1,16'h0045,16'h0189,-16'h0144,16'h0084,16'h0023,-16'h0027,16'h0184,-16'h00cb,16'h01a7,-16'h003b,16'h0113,16'h00c8,-16'h0094,16'h010a,-16'h0016,16'h00cf,-16'h0071,-16'h0082,-16'h001c,-16'h005c,16'h00a4,16'h0002,-16'h0022,-16'h006b,16'h0025,-16'h002c,-16'h004f,-16'h00b8,16'h0017,-16'h001a,-16'h0073,-16'h00db,16'h0067,16'h003c,16'h0109,-16'h019e,16'h002d,16'h012f,16'h0143,-16'h00c3,16'h0028,16'h00ab,-16'h00c0,16'h0058,16'h0135,-16'h00f7,-16'h00ad,-16'h002e,16'h000e,16'h0033,16'h010b,16'h0157,16'h005d,16'h008d,-16'h00c8,-16'h0059,16'h007c,16'h0056,16'h0195,-16'h0084,-16'h00bc,-16'h00c1,16'h0021,-16'h012b,16'h0062,16'h0136,-16'h0109,16'h0000,16'h0054,-16'h0166,16'h0126,-16'h0073,16'h01c6,-16'h0067,16'h014c,16'h0057,-16'h00a4,16'h01da,16'h0054,16'h00bc,-16'h0219,-16'h00d1,-16'h006d,16'h005a,16'h00cb,16'h0006,-16'h0055,-16'h006f,16'h0028,16'h003f,16'h0007,-16'h008f,16'h003f,-16'h0042,-16'h0028,-16'h010a,-16'h0026,-16'h0087,16'h0193,-16'h014a,16'h0024,16'h00f6,16'h00a6,-16'h0102,-16'h007d,16'h0070,-16'h0007,16'h00b3,16'h00ed,-16'h015e,-16'h0056,16'h000e,16'h0058,16'h008a,16'h014d,16'h0139,16'h0073,16'h00a4,-16'h00de,-16'h00d3,16'h0010,-16'h014a,16'h0178,-16'h0039,-16'h0024,-16'h005c,-16'h0011,-16'h0192,16'h00f5,16'h0128,-16'h0063,16'h00ab,16'h0090,-16'h0125,16'h0121,-16'h0051,16'h010f,-16'h00ae,16'h0123,16'h0068,-16'h009a,16'h01a1,16'h0133,16'h00b2,-16'h0222,-16'h0179,-16'h0035,16'h0059,16'h00f8,-16'h0053,-16'h003e,16'h001d,16'h0064,16'h002d,16'h000a,-16'h0112,-16'h0056,-16'h0093,-16'h00c4,-16'h0101,16'h0003,-16'h001a,16'h015d,-16'h0083,16'h0039,16'h00f6,16'h0113,-16'h0186,16'h000d,16'h00ae,16'h0131,16'h00df,16'h00e0,-16'h010b,-16'h00ee,16'h0020,16'h007d,16'h010d,16'h011c,16'h016f,16'h00bc,16'h0067,-16'h001d,-16'h0093,16'h0035,-16'h0186,16'h00ef,-16'h001f,-16'h0063,16'h000c,-16'h002b,-16'h0118,16'h0068,16'h0169,16'h00af,16'h0062,-16'h0009,-16'h00c8,16'h01aa,-16'h002d,16'h0083,-16'h009a,16'h0160,16'h00eb,-16'h005a,16'h019d,16'h00b7,16'h00a2,-16'h01d6,-16'h0278,-16'h0067,16'h0005,16'h0182,16'h0021,-16'h007a,16'h0047,-16'h003e,16'h006e,16'h007b,-16'h00d6,16'h003e,-16'h0086,-16'h005e,-16'h00bb,-16'h0010,-16'h002b,16'h010d,-16'h0079,-16'h0026,-16'h0014,16'h00f1,-16'h01c5,-16'h0011,16'h009e,16'h0109,16'h0148,16'h00d3,-16'h0172,-16'h00dd,-16'h007c,16'h0081,16'h0116,16'h0165,16'h0144,16'h006d,16'h0013,-16'h0012,-16'h00c6,-16'h0009,-16'h01eb,16'h00e4,16'h00bf,-16'h001f,-16'h0034,16'h0055,-16'h011e,-16'h0043,16'h014d,16'h017e,-16'h0028,-16'h0058,-16'h005b,16'h01aa,-16'h0026,-16'h0107,-16'h00ac,16'h013f,16'h0076,-16'h0061,16'h019f,16'h0026,16'h0075,-16'h012e,-16'h02b2,16'h0016,-16'h0029,16'h01a7,16'h0053,16'h000e,-16'h00a7,16'h003d,16'h019c,16'h00a1,-16'h008c,16'h000a,-16'h0077,-16'h004c,-16'h0057,16'h0063,-16'h001f,16'h00dd,16'h0009,-16'h0097,-16'h009b,16'h00da,-16'h0202,16'h0011,16'h00db,16'h01b2,16'h00fa,16'h014c,-16'h0142,-16'h015e,16'h0014,-16'h002e,16'h0044,16'h0124,16'h0133,-16'h001d,-16'h0042,-16'h0015,-16'h0109,-16'h002c,-16'h00f5,16'h0108,16'h0096,-16'h0075,-16'h000d,16'h0049,-16'h0106,-16'h0001,16'h014f,16'h01c3,-16'h00bd,-16'h00d5,16'h0010,16'h01d9,16'h0092,-16'h0293,-16'h0054,16'h0138,16'h0091,-16'h0071,16'h0180,-16'h0068,-16'h004e,-16'h01b8,-16'h00f0,16'h0015,16'h000b,16'h0232,16'h0030,-16'h007d,-16'h0089,16'h0006,16'h010c,-16'h0068,-16'h002c,-16'h002d,16'h00dd,-16'h00f0,-16'h0088,-16'h0004,-16'h00cd,16'h007f,-16'h004d,-16'h0051,-16'h01a4,16'h00fb,-16'h0225,16'h0019,16'h00f6,16'h020d,16'h014b,16'h0136,-16'h00cc,-16'h0254,16'h0122,16'h0015,16'h0056,-16'h0076,16'h00ba,16'h0009,-16'h004a,-16'h0021,-16'h007f,-16'h0095,-16'h0011,16'h0096,16'h0023,-16'h01dc,-16'h00df,16'h0053,-16'h011a,16'h0025,16'h00d0,16'h0106,-16'h004a,-16'h00aa,16'h0003,16'h00f4,16'h008b,-16'h011e,-16'h00c9,16'h01b4,16'h0045,-16'h0069,16'h014a,-16'h0022,-16'h0067,-16'h0187,16'h00d2,16'h0094,-16'h00b5,16'h0248,-16'h000e,-16'h003c,-16'h0072,16'h009a,16'h0133,-16'h002e,-16'h0032,-16'h002d,16'h0224,-16'h00d0,-16'h00b4,16'h004e,-16'h013e,-16'h0051,-16'h009f,16'h0030,-16'h01ce,16'h00c1,-16'h01fb,16'h0077,16'h006e,16'h021c,-16'h0018,16'h0147,-16'h0197,-16'h0314,16'h00d8,16'h004e,-16'h00a2,-16'h01b6,16'h0065,16'h0046,16'h0071,-16'h004a,-16'h000e,-16'h007a,16'h00a5,16'h009b,16'h002d,-16'h01a3,-16'h0047,16'h0041,-16'h00d4,-16'h005d,16'h00e6,16'h010e,-16'h00b0,-16'h008a,-16'h002b,16'h002f,16'h00bb,16'h0189,-16'h0069,16'h0115,16'h0033,16'h0072,16'h00d9,16'h0035,-16'h00a7,-16'h00f9,16'h00e3,-16'h0058,-16'h0140,16'h022b,-16'h00f3,-16'h000d,-16'h008c,16'h00e7,16'h019b,-16'h012e,-16'h0038,16'h003a,16'h011a,-16'h016f,-16'h00e2,16'h001f,-16'h0097,-16'h0057,-16'h0043,16'h0075,-16'h00de,16'h0036,-16'h0121,16'h0099,16'h010a,16'h021f,-16'h016c,16'h011c,-16'h0132,-16'h03e8,16'h007e,16'h00db,-16'h006c,-16'h01b8,16'h0039,-16'h0059,-16'h004e,-16'h0015,16'h0012,-16'h0091,16'h016d,16'h001f,-16'h0038,-16'h0166,-16'h002f,16'h0101,-16'h009b,-16'h008b,16'h0098,16'h003f,-16'h0022,-16'h006a,-16'h0043,-16'h00d2,16'h00cd,16'h02ab,-16'h001d,16'h0144,16'h003c,16'h000d,16'h00d7,16'h007f,-16'h008d,-16'h007b,16'h0148,-16'h006d,-16'h0103,16'h015b,-16'h00f7,-16'h002d,-16'h0098,16'h00c2,16'h0154,-16'h02e2,-16'h00e2,16'h000c,-16'h016d,-16'h0101,-16'h0097,16'h0093,-16'h00c6,16'h005c,16'h004c,16'h0143,-16'h008f,16'h006e,-16'h0032,16'h00fd,16'h0152,16'h0289,-16'h0157,16'h015f,-16'h00af,-16'h043b,16'h00a9,16'h009f,-16'h012d,-16'h0031,16'h0032,-16'h0064,16'h00a6,16'h0041,16'h0078,-16'h0068,16'h00ed,-16'h00ab,-16'h0056,-16'h0128,-16'h0010,16'h00ff,-16'h00a4,-16'h0076,16'h007b,16'h0030,-16'h0014,-16'h0100,-16'h0080,-16'h011a,16'h00e7,16'h01ee,-16'h0088,16'h00fe,16'h001c,16'h0034,16'h00ca,16'h001b,-16'h00aa,16'h00cb,16'h013d,-16'h009a,16'h0051,16'h0180,-16'h00d0,-16'h0072,-16'h00a6,16'h00a3,16'h015b,-16'h03a1,-16'h00c5,16'h00a5,-16'h02f8,16'h00c1,-16'h00e6,16'h0076,-16'h00d3,-16'h002a,16'h002a,16'h0136,-16'h0023,16'h0042,-16'h0032,16'h0164,16'h013e,16'h01c3,-16'h002f,16'h019d,16'h0011,-16'h0423,16'h00aa,16'h005b,-16'h0071,16'h00cf,16'h0008,-16'h00cf,16'h0113,16'h0036,16'h0089,-16'h0078,16'h0130,-16'h00a9,-16'h00d8,-16'h012d,16'h0026,16'h00fe,-16'h0078,-16'h0069,16'h00a1,16'h0066,16'h001d,-16'h0023,-16'h0127,-16'h0011,16'h00c5,16'h00af,-16'h00b5,16'h00cf,16'h0095,16'h0069,16'h00a7,16'h0097,-16'h000a,16'h00ff,16'h0106,-16'h008d,16'h010e,16'h01a9,-16'h00cb,-16'h003f,-16'h001d,16'h0052,16'h0230,-16'h01a4,-16'h0090,16'h002f,-16'h02d2,16'h01a7,-16'h00bc,-16'h0063,-16'h00ee,-16'h000f,16'h0023,16'h01a0,16'h004f,-16'h0055,16'h0074,16'h013c,16'h01f9,16'h01f4,-16'h0075,16'h01a8,16'h001e,-16'h037a,16'h013f,16'h0037,-16'h0050,16'h014d,-16'h0006,-16'h00b6,16'h00e8,16'h006a,16'h00d9,-16'h004c,16'h0114,-16'h00b8,-16'h0115,-16'h00ec,16'h0057,16'h00d0,-16'h0018,-16'h00b7,16'h004d,16'h00a6,16'h008b,16'h0086,-16'h012a,-16'h00b1,16'h0051,-16'h00e1,-16'h00bc,16'h00a2,-16'h0081,16'h0021,16'h00b1,16'h006b,16'h00f4,16'h0102,16'h007b,-16'h006b,16'h0176,16'h0174,-16'h002f,-16'h00c8,16'h010e,-16'h001e,16'h0107,-16'h00b3,-16'h00b4,16'h0066,-16'h0122,16'h01cb,-16'h009d,-16'h0081,-16'h0094,16'h002b,-16'h0083,16'h00d7,16'h0013,-16'h00ea,16'h0085,16'h00c7,16'h0155,16'h0130,-16'h0022,16'h01ec,16'h0082,-16'h0336,16'h01a8,16'h008c,-16'h0060,16'h01ec,16'h0047,-16'h005b,16'h00f1,16'h0003,16'h0103,-16'h00d9,16'h00d6,-16'h00ab,-16'h00f0,-16'h0114,16'h0028,16'h010d,-16'h00bd,-16'h008d,16'h00c2,-16'h0083,16'h0081,16'h019a,-16'h0061,-16'h0111,16'h0001,-16'h022e,-16'h011f,16'h0090,-16'h008f,-16'h002a,16'h0056,16'h006a,16'h015c,16'h010a,16'h0009,-16'h0012,16'h022a,16'h0207,-16'h000c,-16'h00a5,16'h00fe,16'h0000,-16'h0024,-16'h0026,-16'h0115,16'h0060,-16'h004b,-16'h009c,-16'h0115,16'h0032,-16'h004b,16'h004b,-16'h00de,-16'h0063,-16'h0019,-16'h004b,-16'h001f,16'h00a0,16'h016e,16'h011a,-16'h00a3,16'h013e,16'h0152,-16'h02f8,16'h0158,16'h0055,16'h000a,16'h01c8,16'h004d,-16'h0024,16'h00e5,16'h0017,16'h00c6,-16'h00b9,16'h00c1,-16'h00e7,-16'h0153,-16'h00e5,16'h0027,16'h011c,-16'h00a1,-16'h0049,16'h0045,-16'h0164,16'h011b,16'h00d8,-16'h0059,-16'h00de,16'h0014,-16'h014e,-16'h0126,16'h003d,-16'h000a,16'h0029,-16'h0009,16'h00ef,16'h0159,16'h0091,-16'h001a,-16'h003e,16'h018d,16'h0205,16'h0088,-16'h0080,16'h0086,16'h001c,-16'h013c,16'h00ae,-16'h0139,-16'h0077,16'h0029,-16'h03aa,-16'h0058,16'h0011,-16'h00ad,-16'h0035,-16'h0060,-16'h00c9,16'h0012,16'h007c,16'h0013,16'h00bd,16'h010a,16'h013b,-16'h0044,16'h011e,16'h00d7,-16'h02c1,16'h012f,16'h00cd,16'h003a,16'h00ca,16'h0101,-16'h001a,16'h001f,16'h0007,16'h00ee,-16'h00ed,16'h0071,16'h0058,-16'h00b7,-16'h006e,16'h002a,16'h017c,-16'h0083,16'h002b,16'h00b2,-16'h0102,16'h007f,16'h0041,-16'h004a,-16'h0078,16'h001b,-16'h0069,-16'h0043,-16'h000a,16'h0033,16'h0044,-16'h0070,16'h00d2,16'h010d,16'h00c3,-16'h015d,-16'h0062,16'h00d3,16'h019d,16'h00a9,-16'h0058,16'h002e,16'h00a3,-16'h0125,16'h0151,-16'h011a,-16'h01b2,16'h00bb,-16'h03e4,16'h004a,16'h00f5,-16'h009e,-16'h001d,-16'h003c,-16'h00cd,-16'h004d,-16'h0051,-16'h0023,16'h0088,16'h0114,16'h0119,-16'h0021,16'h00ef,16'h00a7,-16'h0247,16'h0156,16'h012a,-16'h00fe,16'h00a5,16'h0091,-16'h000e,-16'h0026,-16'h001e,16'h00dd,-16'h00fb,16'h001b,-16'h0026,-16'h0074,-16'h00ea,16'h0051,16'h012e,-16'h008a,16'h0140,16'h00e0,-16'h0136,16'h00d8,16'h0084,16'h0037,16'h0085,-16'h0081,16'h01a0,16'h008b,-16'h0011,16'h0043,-16'h0013,-16'h003e,16'h00be,16'h004e,16'h0091,-16'h024b,-16'h0034,-16'h0039,16'h01ab,16'h0165,-16'h00d1,-16'h0089,16'h007e,-16'h0189,16'h00e6,-16'h012a,-16'h0214,16'h00b3,-16'h01cd,16'h005b,16'h008a,-16'h00db,16'h004e,-16'h0010,-16'h0039,-16'h00e3,-16'h0039,-16'h0051,16'h00d6,16'h0050,16'h014a,16'h00ae,16'h003a,16'h006d,-16'h01ab,16'h0118,16'h01e0,-16'h00d6,-16'h00a6,16'h008a,-16'h00fe,-16'h0051,16'h003f,16'h00d8,-16'h012e,-16'h0074,16'h0004,16'h0000,-16'h0159,-16'h0020,16'h00f7,-16'h0029,16'h0123,16'h00b0,-16'h00ff,16'h00d7,16'h00f8,16'h00dc,16'h0057,-16'h00a6,16'h014f,16'h0132,16'h005c,16'h0090,16'h0015,-16'h0052,16'h006f,-16'h00d5,16'h00ca,-16'h0270,-16'h0056,-16'h00a3,16'h014e,16'h0163,-16'h0077,-16'h0068,16'h0041,-16'h015b,16'h008f,-16'h015d,-16'h01d2,-16'h0044,16'h0161,16'h001d,16'h00da,-16'h00f5,16'h013d,16'h002f,-16'h0105,-16'h0110,-16'h000e,-16'h0082,16'h003c,16'h0045,16'h00e9,16'h00cb,16'h0026,16'h009f,-16'h0174,16'h0117,16'h023f,-16'h00a4,-16'h0163,16'h008d,-16'h00fa,16'h004d,-16'h0042,-16'h002a,-16'h0115,-16'h005d,16'h005d,-16'h0004,-16'h01d8,16'h001e,16'h00e1,16'h002d,16'h00aa,16'h006a,-16'h001a,16'h00cf,16'h0043,16'h00e8,16'h0009,-16'h0073,16'h0119,16'h01e9,16'h0031,16'h0098,16'h0046,-16'h001d,16'h0138,-16'h0181,-16'h002e,-16'h015c,-16'h006b,-16'h006a,16'h012f,16'h0116,-16'h00cc,-16'h00b8,16'h004a,-16'h00fe,-16'h0026,-16'h00f5,-16'h00a0,16'h0019,16'h018b,16'h0055,-16'h00b4,-16'h0131,16'h011a,16'h0036,-16'h010a,-16'h019f,16'h0001,-16'h013d,-16'h0074,-16'h0057,16'h009e,16'h010d,-16'h0001,-16'h003a,-16'h0148,16'h00a6,16'h0227,16'h00bf,-16'h00e9,16'h00b7,-16'h0126,16'h00c1,-16'h0098,-16'h0041,-16'h011a,16'h0052,16'h006b,16'h0104,-16'h0158,16'h0015,16'h00c5,16'h0000,16'h0076,16'h00b2,16'h0063,16'h00a7,-16'h000e,16'h009c,16'h0075,-16'h0074,16'h00da,16'h0181,16'h0019,16'h0068,16'h008a,16'h0011,16'h00b5,-16'h03d8,-16'h0016,-16'h0109,-16'h0034,-16'h008e,16'h00c7,16'h007d,-16'h013e,-16'h0072,16'h00ba,-16'h0017,-16'h009f,-16'h010a,16'h00a8,-16'h0016,16'h0138,16'h00c3,-16'h0244,-16'h00ee,16'h0120,-16'h0082,-16'h0014,-16'h01d8,-16'h0099,-16'h018a,-16'h0082,-16'h0066,16'h002b,16'h0133,-16'h0078,-16'h0057,-16'h0142,-16'h006d,16'h0129,16'h00fb,-16'h0073,16'h00e7,-16'h00f9,16'h0162,-16'h0073,-16'h008c,-16'h00e6,16'h004d,16'h0097,-16'h000d,-16'h01ac,16'h0046,16'h0121,16'h0035,16'h0056,16'h00a9,16'h0056,16'h00f8,16'h0069,16'h0087,16'h0065,-16'h009c,16'h0054,-16'h0073,-16'h0103,-16'h001a,16'h0086,16'h0076,16'h0013,-16'h0588,-16'h007c,-16'h00a2,-16'h002a,16'h0021,16'h00c9,16'h0042,-16'h0138,16'h009c,16'h00df,16'h0032,-16'h0174,-16'h0049,16'h01b8,16'h0054,16'h01b6,16'h0040,-16'h0245,-16'h00d7,16'h007a,-16'h00a4,16'h0110,-16'h01ba,-16'h00db,-16'h01a1,16'h0007,-16'h001e,-16'h0078,16'h01d5,-16'h0048,-16'h0053,-16'h00f9,16'h0007,16'h0052,16'h0107,-16'h002d,16'h0119,-16'h0054,16'h01d2,-16'h0013,-16'h001c,-16'h011b,-16'h003b,16'h0011,-16'h0140,-16'h0203,16'h00d3,16'h00fe,-16'h0067,16'h00a9,16'h011f,16'h0061,16'h00dd,16'h00bc,-16'h0007,16'h0055,-16'h009e,16'h0086,-16'h034e,-16'h0121,-16'h00f5,16'h0075,16'h005f,-16'h002b,-16'h0420,-16'h00be,-16'h006b,-16'h0011,16'h0057,16'h0137,-16'h005b,-16'h00dd,16'h0114,16'h00b3,16'h0039,-16'h00e3,-16'h0025,16'h018b,16'h0079,-16'h0034,16'h0010,-16'h018e,-16'h00be,16'h0062,-16'h0055,16'h0147,-16'h00aa,16'h002c,-16'h0188,16'h0050,-16'h006c,-16'h002d,16'h00fb,16'h0045,-16'h013e,-16'h00e3,16'h0061,-16'h01e8,16'h0161,-16'h004c,16'h00dc,-16'h006d,16'h0233,16'h0087,16'h0065,-16'h0113,16'h003c,-16'h0021,-16'h02be,-16'h0237,16'h01db,16'h005b,-16'h00df,16'h012d,16'h011a,16'h00ad,16'h011e,16'h004d,16'h0094,-16'h0053,-16'h00f1,16'h0022,-16'h05c2,-16'h0110,-16'h0147,16'h008a,16'h00be,-16'h00ce,-16'h0282,-16'h0024,-16'h0047,-16'h0033,16'h0028,16'h014f,-16'h0137,-16'h0083,16'h00ff,16'h0017,16'h0031,-16'h0065,-16'h008a,16'h00af,16'h00b3,-16'h02a2,16'h0023,16'h005a,-16'h00b0,16'h004c,-16'h000d,16'h0128,-16'h003b,-16'h0035,-16'h014c,-16'h006f,16'h0050,-16'h0010,16'h00a0,16'h0088,-16'h00df,-16'h0022,-16'h005a,-16'h02ab,16'h01b3,-16'h0005,16'h009d,-16'h0004,16'h00c8,16'h0092,16'h00df,-16'h0103,-16'h005c,16'h009a,-16'h03d8,-16'h0262,16'h01c1,16'h0091,-16'h00b8,16'h01eb,16'h0209,16'h000d,16'h00ea,16'h0077,-16'h0082,-16'h0004,-16'h008a,-16'h000b,-16'h0574,-16'h00d8,-16'h008d,16'h0003,16'h013f,-16'h00a8,-16'h01cb,-16'h0054,-16'h0076,-16'h0082,16'h001d,16'h01b4,-16'h02b4,-16'h0078,16'h0065,-16'h0015,-16'h0058,-16'h0059,-16'h0068,-16'h00ab,-16'h0004,-16'h02b1,16'h0032,16'h01dd,-16'h008a,16'h0026,16'h0098,16'h018a,-16'h0014,-16'h014c,-16'h01a4,-16'h0041,16'h0045,16'h0092,-16'h000f,16'h00d4,-16'h0085,-16'h0096,-16'h00e0,-16'h019b,16'h01f1,16'h0024,16'h00a0,-16'h008a,-16'h0034,16'h002a,16'h00aa,-16'h00e5,16'h000f,16'h007e,-16'h02b6,-16'h033b,16'h0233,-16'h0001,-16'h0055,16'h013b,16'h01e4,-16'h0085,16'h0116,16'h00c9,-16'h0080,16'h00b0,16'h0019,16'h0015,-16'h03c6,-16'h0094,-16'h0034,-16'h0128,16'h00d6,-16'h0037,-16'h012b,-16'h009f,-16'h00ea,-16'h00c8,16'h0028,16'h0135,-16'h040c,16'h000a,-16'h0071,-16'h0146,-16'h0082,-16'h0023,-16'h0145,-16'h01ee,16'h0060,-16'h00d1,-16'h0003,16'h02d9,-16'h0059,-16'h00a7,16'h0015,16'h015e,-16'h0033,-16'h0209,-16'h01bd,-16'h002c,-16'h000b,-16'h0015,-16'h001b,16'h0130,16'h000d,-16'h007a,-16'h00e5,-16'h0128,16'h0125,16'h004d,16'h00f1,-16'h00b7,-16'h020e,16'h0050,16'h0030,-16'h00f7,-16'h000d,16'h0017,-16'h027f,-16'h0340,16'h018c,-16'h001b,-16'h0099,16'h00aa,16'h0104,-16'h014f,16'h0108,16'h00a9,-16'h0021,16'h005e,16'h0067,16'h000c,-16'h006a,-16'h00a0,16'h0124,-16'h014d,16'h00a0,16'h0031,-16'h00e8,-16'h00e6,-16'h0061,16'h002f,16'h0057,16'h018a,-16'h036e,16'h000a,-16'h0120,-16'h03f2,-16'h0018,-16'h0037,-16'h0173,-16'h02c8,16'h0027,16'h010c,16'h0103,16'h0240,16'h0040,-16'h00ff,16'h0026,16'h0187,16'h0029,-16'h0124,-16'h01b2,16'h001b,16'h005c,-16'h0002,16'h006f,16'h015d,-16'h004e,16'h0009,-16'h00fc,-16'h0032,16'h0167,16'h003d,16'h0094,-16'h00f6,-16'h02e0,-16'h0024,-16'h0014,-16'h0054,16'h001e,16'h0127,-16'h01de,-16'h031e,16'h00fb,16'h0019,-16'h011c,16'h011f,16'h0162,-16'h00df,16'h00ef,16'h0155,-16'h00aa,16'h004f,16'h008e,-16'h00f3,16'h01a6,-16'h0120,16'h0223,-16'h011a,-16'h0073,16'h0090,-16'h00ce,-16'h0179,-16'h0126,16'h0051,16'h00bb,16'h0116,-16'h01a4,-16'h005f,-16'h00f4,-16'h04b6,16'h004d,-16'h0052,-16'h0293,-16'h0297,-16'h0018,16'h00ee,16'h0229,16'h0084,-16'h0023,-16'h015c,16'h01ac,16'h01c0,16'h0196,-16'h012f,-16'h018c,16'h008e,16'h012e,-16'h000e,16'h00ba,16'h0128,-16'h0071,16'h0058,16'h0000,-16'h011e,16'h01b3,16'h0011,16'h00df,-16'h00bc,-16'h0176,-16'h00c4,-16'h00b3,-16'h004d,16'h009e,16'h00fc,-16'h016e,-16'h036c,-16'h0044,-16'h0028,-16'h0188,16'h00b1,16'h0156,-16'h0059,16'h017f,16'h00dd,-16'h0104,16'h013b,16'h001f,-16'h0072,16'h02c3,-16'h0160,16'h0191,-16'h00fd,-16'h0099,16'h0177,16'h0001,-16'h0176,-16'h0113,16'h0115,-16'h000e,16'h00ed,-16'h0024,-16'h00ec,-16'h0076,-16'h02d7,16'h00d5,-16'h0034,-16'h033b,-16'h0180,16'h0053,16'h0133,16'h02b7,-16'h0036,-16'h0091,-16'h01b1,16'h01d4,16'h0254,16'h0180,-16'h0118,-16'h019a,16'h007b,16'h0215,16'h009f,16'h00b2,16'h00b6,-16'h0140,-16'h004f,-16'h003e,-16'h0169,16'h00e2,16'h0029,16'h0194,-16'h00db,-16'h0065,16'h0056,-16'h0164,-16'h00a6,-16'h0043,16'h0190,-16'h0108,-16'h0015,-16'h0139,-16'h00e5,-16'h013a,-16'h003e,16'h01c9,-16'h0070,-16'h001e,-16'h001e,16'h0056,16'h026d,-16'h0093,16'h00f7,16'h007e,16'h00d9,16'h0024,-16'h0045,-16'h0034,16'h000b,16'h00db,-16'h0007,-16'h0030,16'h0008,-16'h006e,16'h0060,-16'h0030,16'h007d,-16'h008e,16'h0018,16'h0089,-16'h005a,-16'h001e,-16'h00b7,16'h00f1,-16'h0016,-16'h0054,16'h0046,-16'h0040,16'h01ea,-16'h00f1,16'h0065,16'h0129,16'h0192,-16'h002a,-16'h00f4,16'h0071,-16'h0124,16'h0014,16'h0160,-16'h0065,-16'h0084,-16'h007d,-16'h00a4,16'h0047,16'h0137,16'h017b,16'h0136,-16'h000e,-16'h00c5,16'h00a0,16'h00fc,-16'h0045,16'h0260,-16'h0043,-16'h0047,-16'h00ca,-16'h00c5,-16'h010c,16'h001d,16'h0141,-16'h00cf,16'h0074,-16'h001b,-16'h009f,16'h021d,-16'h005e,16'h0129,16'h0006,16'h0104,16'h00a1,-16'h00d0,16'h00b3,16'h0056,16'h005d,-16'h0065,-16'h0114,-16'h003e,-16'h0004,16'h0029,-16'h0047,-16'h0031,-16'h0081,-16'h001c,16'h000f,-16'h0008,-16'h0023,16'h0002,16'h0020,16'h0008,-16'h0100,16'h0012,16'h002c,16'h0186,-16'h0173,-16'h0028,16'h016f,16'h0141,-16'h00ce,16'h0027,16'h00af,-16'h00a6,16'h004d,16'h00f3,-16'h0077,16'h003c,-16'h006f,16'h006f,-16'h006a,16'h014a,16'h019c,16'h0082,16'h004c,-16'h0092,-16'h0003,16'h011d,-16'h0037,16'h0202,16'h000f,-16'h002d,-16'h0074,-16'h012d,-16'h0141,16'h0092,16'h00fc,-16'h0097,16'h008c,-16'h000a,-16'h0182,16'h01f4,-16'h0066,16'h0148,-16'h0095,16'h0167,16'h0057,-16'h00a4,16'h015d,16'h0059,16'h0088,-16'h0181,-16'h011d,-16'h007b,16'h0007,16'h0062,-16'h007e,-16'h0041,-16'h0093,16'h0031,16'h0090,16'h0088,-16'h0032,16'h005c,-16'h0078,16'h0009,-16'h009a,-16'h0017,-16'h00b1,16'h0131,-16'h0164,16'h000d,16'h0145,16'h014c,-16'h005c,-16'h005b,16'h010f,16'h0004,16'h007b,16'h00e6,-16'h011d,-16'h003e,-16'h0045,16'h0025,16'h00ce,16'h019b,16'h016a,16'h0075,16'h00ad,-16'h0041,16'h0019,16'h00b3,-16'h012d,16'h0159,-16'h0011,16'h0020,-16'h0099,-16'h01a6,-16'h00ee,16'h0095,16'h01a7,16'h0018,16'h006f,-16'h0034,-16'h01a7,16'h017b,-16'h0007,16'h00b9,-16'h0083,16'h0100,16'h0135,-16'h0053,16'h022a,16'h0154,16'h00c9,-16'h0218,-16'h0190,-16'h005e,16'h008e,16'h0091,-16'h0038,-16'h0089,-16'h001d,-16'h0029,16'h0043,16'h00e6,-16'h00f0,16'h007f,-16'h00ef,-16'h002d,-16'h0199,-16'h0074,-16'h00ad,16'h0198,-16'h002c,16'h000e,16'h001e,16'h010c,-16'h0094,-16'h0006,16'h0044,16'h00de,16'h0082,16'h0101,-16'h0081,-16'h004e,16'h0020,16'h0045,16'h0081,16'h0141,16'h01d1,16'h00fe,16'h00e2,-16'h0021,-16'h0027,16'h005e,-16'h0164,16'h016a,16'h0018,-16'h001d,-16'h0023,-16'h01a4,-16'h0187,16'h004f,16'h0176,16'h0030,16'h007e,-16'h0011,-16'h0127,16'h028f,-16'h001a,16'h0000,-16'h005f,16'h0167,16'h0130,16'h0016,16'h02b3,16'h00dc,16'h0088,-16'h0262,-16'h0286,-16'h0055,-16'h0058,16'h014b,16'h004e,-16'h002d,-16'h0011,-16'h0067,16'h00b6,16'h0098,-16'h00b9,16'h005d,-16'h00f9,-16'h008c,-16'h00e9,-16'h0039,-16'h008b,16'h015a,16'h0044,16'h0029,-16'h0080,16'h00eb,-16'h0059,16'h0038,16'h0072,16'h00d5,16'h009e,16'h00d2,-16'h0169,-16'h00d5,16'h0005,-16'h001e,16'h002d,16'h0164,16'h0103,16'h00d8,16'h0032,-16'h0069,16'h0003,16'h0053,-16'h012d,16'h0156,16'h00d2,16'h003f,16'h0023,-16'h01d7,-16'h00ea,16'h0032,16'h0148,16'h0102,-16'h0022,-16'h00ba,-16'h00ba,16'h0211,-16'h002c,-16'h01c0,-16'h005d,16'h0123,16'h0132,-16'h0021,16'h0206,-16'h0016,-16'h0004,-16'h0186,-16'h01c1,-16'h0017,-16'h00cd,16'h016d,-16'h000d,-16'h0036,16'h0005,-16'h0092,16'h010c,-16'h0015,-16'h00d2,-16'h0001,16'h0011,16'h003b,-16'h0099,-16'h0048,-16'h0085,16'h00d8,-16'h0075,16'h008e,-16'h0136,16'h0095,-16'h000e,-16'h004e,16'h0081,16'h00b8,16'h0029,16'h0142,-16'h00a3,-16'h010f,16'h0054,-16'h0006,-16'h0064,16'h00b1,16'h0049,-16'h000d,-16'h0009,-16'h001e,16'h0030,-16'h000d,-16'h0010,16'h0124,16'h006c,-16'h0050,16'h0046,-16'h0156,-16'h0108,16'h00b6,16'h010f,16'h00c0,-16'h0092,-16'h00b3,-16'h0075,16'h01d5,16'h005a,-16'h0175,-16'h0039,16'h0135,16'h00eb,16'h0005,16'h0252,16'h000f,-16'h0015,-16'h0125,-16'h0006,16'h0028,-16'h0091,16'h0191,-16'h0041,-16'h0073,16'h0029,16'h000f,16'h0123,16'h0006,-16'h00a5,-16'h009c,16'h012a,-16'h00bd,-16'h00aa,-16'h0004,-16'h00a4,16'h0081,-16'h0078,16'h0021,-16'h0223,16'h0156,-16'h006a,16'h001b,16'h012d,16'h00b0,16'h0126,16'h01a2,-16'h0118,-16'h0172,16'h00bf,16'h004a,-16'h00d4,-16'h00bc,16'h0097,16'h001b,16'h0033,16'h0004,16'h002b,-16'h0036,16'h00db,16'h009d,16'h0038,-16'h015b,-16'h0078,-16'h01c4,-16'h011d,16'h0087,16'h00e9,16'h00a6,-16'h0033,-16'h0063,-16'h0048,16'h0048,16'h00a5,-16'h0027,16'h002a,16'h012a,16'h0087,16'h003d,16'h027b,-16'h000c,-16'h003f,-16'h0125,16'h0101,-16'h004c,-16'h00fb,16'h00a2,-16'h008d,-16'h0020,16'h004b,16'h00bb,16'h00eb,-16'h019f,-16'h009b,-16'h0041,16'h01d3,-16'h00bb,-16'h00c2,-16'h002e,-16'h0116,16'h0000,-16'h004c,16'h0078,-16'h0221,16'h00a6,-16'h007f,-16'h001d,16'h00c6,16'h00f0,16'h0060,16'h0183,-16'h00b7,-16'h011a,16'h00a6,-16'h0010,-16'h0168,-16'h0161,16'h000d,16'h00b5,16'h00ce,-16'h0003,16'h0058,16'h0011,16'h013c,16'h00e5,16'h0033,-16'h0185,-16'h00ec,-16'h015f,-16'h0172,-16'h0003,16'h0060,16'h004f,-16'h0011,-16'h0035,-16'h00c5,16'h0046,16'h0061,16'h01f0,16'h000d,16'h00ed,16'h008b,16'h0057,16'h0185,16'h002f,-16'h00a3,-16'h0074,16'h0092,-16'h014c,-16'h00f4,16'h0099,-16'h011d,-16'h0074,-16'h0086,16'h0086,16'h00ed,-16'h02d8,-16'h013d,16'h0040,16'h0072,-16'h012a,-16'h006b,16'h0000,-16'h00cc,16'h0039,-16'h0080,16'h014a,-16'h01c3,16'h0033,-16'h004a,-16'h003c,16'h014c,16'h011e,-16'h00e9,16'h0125,-16'h010a,-16'h0166,16'h0062,16'h007c,-16'h01ec,-16'h0185,16'h0046,-16'h000d,16'h00ab,16'h0041,16'h002c,16'h0041,16'h0184,16'h006a,-16'h002b,-16'h01e5,-16'h010d,-16'h0088,-16'h0161,-16'h0080,16'h00a7,-16'h0041,-16'h0042,-16'h00b7,-16'h01c5,-16'h0076,16'h00e6,16'h0284,16'h0097,16'h00ac,16'h008a,16'h006a,16'h01ee,16'h008a,-16'h0097,16'h0034,16'h011f,-16'h016e,16'h0055,16'h00ce,-16'h018f,-16'h00f5,-16'h0076,16'h0055,16'h00f5,-16'h038e,-16'h0158,16'h007e,-16'h01ee,-16'h009a,-16'h00a9,16'h0044,-16'h0101,-16'h007b,16'h0067,16'h0144,-16'h00ec,16'h00c5,-16'h00ce,16'h00b6,16'h01ac,16'h00f4,-16'h00d7,16'h019f,-16'h000f,-16'h0179,16'h000f,16'h0003,-16'h01d8,16'h0052,-16'h0049,-16'h005e,16'h011b,16'h0066,16'h000c,-16'h005a,16'h0123,-16'h0088,-16'h006b,-16'h00fc,-16'h0061,-16'h0019,-16'h0129,-16'h0022,16'h00ef,-16'h0028,-16'h002d,-16'h0070,-16'h01f1,-16'h0107,16'h0077,16'h0192,-16'h005a,16'h0093,16'h00c9,16'h0043,16'h0245,16'h0095,-16'h010e,16'h0156,16'h00d8,-16'h0117,16'h014d,16'h00bf,-16'h012a,-16'h0052,-16'h0070,16'h0006,16'h015d,-16'h0250,-16'h0164,16'h00db,-16'h031f,16'h0084,-16'h0088,16'h006a,-16'h015e,-16'h0022,-16'h0004,16'h00f1,16'h0034,16'h000c,-16'h006d,16'h0093,16'h01af,16'h006a,-16'h00a2,16'h0195,16'h002f,-16'h0121,16'h003a,-16'h001e,-16'h00f2,16'h0106,-16'h0068,-16'h0060,16'h0108,16'h008b,16'h00bb,-16'h0030,16'h0142,-16'h00d5,-16'h00e8,-16'h00e4,-16'h00da,-16'h0010,-16'h0135,-16'h009e,16'h0077,16'h0064,16'h0001,16'h007e,-16'h01f1,-16'h0116,16'h0044,16'h0023,-16'h0102,16'h0013,16'h0060,16'h002d,16'h01cb,16'h0092,-16'h0046,16'h0111,16'h0074,-16'h013c,16'h022f,16'h00b3,-16'h006a,-16'h0081,16'h005a,-16'h003b,16'h016e,-16'h012a,-16'h01b9,16'h00c7,-16'h02dc,16'h018f,-16'h0066,-16'h0040,-16'h0145,-16'h0034,-16'h000b,16'h00ae,16'h00af,-16'h0053,16'h0028,16'h0120,16'h01e4,16'h00c6,-16'h0079,16'h01b8,16'h0057,-16'h018c,16'h00d7,16'h001e,-16'h0119,16'h0151,16'h004b,-16'h003b,16'h00e8,16'h0071,16'h0109,16'h0018,16'h00e3,-16'h0081,-16'h0064,-16'h014d,-16'h00ab,16'h0008,-16'h01df,-16'h005f,16'h0056,16'h0045,16'h0089,16'h00cc,-16'h0177,-16'h00ea,16'h0069,-16'h016b,-16'h017b,16'h0025,-16'h0048,16'h0012,16'h01b5,16'h006f,16'h0097,16'h011f,16'h0012,-16'h00c8,16'h022f,16'h008e,-16'h001b,-16'h00fb,16'h010f,-16'h0105,16'h005e,-16'h0086,-16'h01a6,16'h0028,-16'h00b0,16'h01e7,-16'h0085,-16'h00c2,-16'h00ea,16'h000f,-16'h00b8,16'h006a,16'h00bc,-16'h004a,16'h0030,16'h0081,16'h016f,-16'h0012,16'h000c,16'h01e1,16'h0146,-16'h0155,16'h00a3,16'h0038,-16'h0133,16'h00f8,-16'h0001,-16'h007a,16'h00db,16'h0068,16'h00a1,-16'h0041,16'h0163,-16'h00a4,-16'h00dd,-16'h00f6,-16'h00db,-16'h0005,-16'h0207,16'h0055,16'h00a1,-16'h010e,16'h00cd,16'h014c,-16'h0155,-16'h00f7,16'h001e,-16'h016f,-16'h0177,-16'h0002,-16'h00c4,-16'h004e,16'h01eb,16'h0063,16'h00f8,16'h00bf,-16'h004e,-16'h00af,16'h0164,16'h00bd,16'h0055,-16'h00b3,16'h015d,-16'h0072,-16'h00c4,16'h0037,-16'h015d,16'h00ca,16'h000f,-16'h0036,-16'h0102,16'h0041,-16'h0159,16'h00c4,-16'h00b3,-16'h0068,16'h003d,16'h0026,-16'h0080,16'h0107,16'h00e4,-16'h0024,-16'h0028,16'h01a5,16'h017f,-16'h018e,16'h0108,16'h005d,-16'h00c7,16'h012d,16'h004b,-16'h0085,16'h006a,-16'h0067,16'h001d,-16'h0090,16'h011a,-16'h0069,-16'h00ce,-16'h0137,-16'h0111,16'h0017,-16'h0232,16'h0029,16'h0095,-16'h00d2,16'h0064,16'h0070,-16'h0170,16'h0016,16'h0047,-16'h0041,-16'h0177,-16'h0021,16'h004b,-16'h0036,16'h0128,16'h0056,16'h00d2,16'h007d,-16'h00d4,-16'h008a,16'h0100,16'h00e9,16'h0056,-16'h00c6,16'h013a,-16'h00b4,-16'h00e7,16'h0040,-16'h01b3,-16'h0060,16'h0008,-16'h0306,-16'h00d4,16'h0116,-16'h00fd,16'h0070,-16'h006d,-16'h00bf,16'h002d,-16'h001c,16'h0037,16'h00eb,16'h0101,-16'h0048,-16'h0010,16'h019b,16'h00ef,-16'h0113,16'h0162,16'h006a,-16'h001c,16'h00b6,16'h003e,16'h006d,16'h007e,-16'h000a,16'h0084,-16'h00ed,16'h01e0,-16'h007a,-16'h00a3,-16'h0126,-16'h005f,-16'h0019,-16'h024e,16'h0057,16'h007f,-16'h00a6,16'h0035,-16'h0007,-16'h0050,16'h00ab,16'h007b,16'h0089,-16'h002b,-16'h0055,16'h003c,-16'h0003,16'h00ce,16'h00ef,16'h0061,16'h00dd,-16'h0112,-16'h00dd,16'h0000,16'h0131,16'h00ae,-16'h00ba,16'h0134,-16'h0020,-16'h0126,16'h0077,-16'h012e,-16'h0216,16'h009b,-16'h032d,-16'h0020,16'h00ab,-16'h0071,16'h009f,-16'h00d6,-16'h017e,16'h0041,16'h0023,16'h002c,16'h0145,16'h0102,-16'h001d,16'h006f,16'h00ef,16'h0049,-16'h016a,16'h0124,16'h016c,-16'h0007,16'h0028,16'h0060,16'h0045,16'h0067,-16'h0095,16'h0034,-16'h014d,16'h015f,16'h003c,16'h0039,-16'h00eb,-16'h0083,-16'h0029,-16'h011a,16'h0181,16'h00d1,-16'h00b6,16'h0095,16'h0020,16'h0030,16'h00e1,16'h0022,16'h0168,16'h00de,16'h0012,16'h0057,-16'h004d,16'h00dc,16'h009b,16'h0028,16'h0086,-16'h00fa,-16'h00e2,-16'h00d7,16'h0132,16'h0045,-16'h013e,16'h003d,16'h000a,-16'h017d,16'h0082,-16'h0158,-16'h031a,16'h0009,-16'h0077,16'h0006,16'h0085,-16'h00a1,-16'h0061,-16'h0066,-16'h00de,-16'h00c0,16'h0072,16'h0081,16'h00d0,16'h007a,-16'h0029,-16'h000a,16'h0092,-16'h001e,-16'h0129,16'h00ec,16'h0188,-16'h001b,-16'h0115,16'h0006,-16'h005d,16'h0062,-16'h0087,-16'h00df,-16'h0152,16'h007f,-16'h0032,16'h00c1,-16'h025a,-16'h0093,-16'h0008,-16'h00d2,16'h0185,16'h009b,-16'h00eb,16'h00a6,16'h0017,16'h0080,16'h0037,16'h0066,16'h0106,16'h0124,-16'h0031,16'h00d4,-16'h003d,16'h00f5,16'h00a8,-16'h0077,16'h0021,-16'h011a,-16'h013c,-16'h008a,16'h00ba,16'h0027,-16'h00e8,-16'h0057,16'h00af,-16'h00f1,16'h005a,-16'h00e0,-16'h02ae,16'h005a,16'h00ac,-16'h0039,16'h003c,-16'h0155,-16'h0010,-16'h0069,-16'h00c4,-16'h0143,-16'h0046,-16'h000b,16'h0053,16'h0035,-16'h0033,16'h00ed,16'h00c4,-16'h0027,-16'h00b4,16'h008f,16'h0203,16'h0059,-16'h00f0,16'h0008,-16'h00e8,16'h0088,-16'h0019,-16'h016c,-16'h00f2,16'h008b,16'h006a,16'h00ec,-16'h01de,-16'h004f,-16'h0044,-16'h00f6,16'h0179,16'h005e,-16'h004d,16'h00a9,16'h0081,16'h00cd,16'h0074,-16'h0008,16'h00e6,16'h016a,16'h0092,16'h00bd,16'h003e,16'h016a,16'h0060,-16'h0124,-16'h004c,-16'h0161,-16'h00c9,-16'h00bf,16'h00b6,16'h005e,-16'h00b6,-16'h0071,16'h00e0,-16'h00cd,16'h0001,-16'h00b4,-16'h017c,16'h0051,16'h0174,-16'h0047,-16'h00d6,-16'h00d7,16'h0054,-16'h0010,-16'h0015,-16'h010e,16'h001c,-16'h00df,-16'h001d,16'h0043,-16'h0069,16'h00a0,16'h0095,16'h0075,-16'h0129,16'h0051,16'h00db,16'h0169,-16'h0119,16'h001a,-16'h0131,16'h009f,-16'h005a,-16'h01f8,-16'h0115,16'h006e,16'h007c,16'h01b2,-16'h01de,-16'h005e,16'h0011,-16'h0081,16'h0130,16'h00e4,16'h004e,16'h00f8,16'h000b,16'h0083,16'h0092,16'h0014,16'h00b6,16'h016d,-16'h0011,16'h00e3,-16'h0047,16'h0150,16'h002c,-16'h0249,-16'h0049,-16'h00a9,-16'h00e5,-16'h00d5,16'h00f4,-16'h0026,-16'h015e,-16'h0016,16'h009a,16'h0054,-16'h004b,-16'h0115,16'h0064,-16'h0055,16'h0196,-16'h0009,-16'h0275,-16'h006e,16'h00aa,-16'h007e,16'h0056,-16'h0146,16'h001d,-16'h01e9,-16'h0050,16'h0024,16'h0012,16'h00db,16'h0005,-16'h0022,-16'h00d5,16'h0002,16'h0031,16'h0192,-16'h004f,16'h0088,-16'h0127,16'h0160,-16'h0004,-16'h01fd,-16'h00ed,-16'h0005,-16'h0066,16'h020b,-16'h02a6,-16'h0065,-16'h0039,-16'h00b9,16'h008b,16'h011d,-16'h0017,16'h00c3,16'h00d3,16'h0093,16'h00a2,-16'h0020,16'h0059,16'h0000,-16'h00a1,16'h0028,-16'h008f,16'h00ef,-16'h00e6,-16'h04ab,-16'h0130,-16'h00b8,-16'h001d,-16'h0021,16'h009e,-16'h0005,-16'h011d,16'h0126,16'h00f4,16'h0084,-16'h0135,-16'h0109,16'h01ab,16'h00d7,16'h0130,16'h003b,-16'h01d4,-16'h00c1,16'h00a8,-16'h00ac,16'h0173,-16'h014c,16'h0058,-16'h0201,16'h007d,16'h0010,-16'h00f3,16'h00d9,16'h0005,16'h0000,-16'h0111,-16'h0058,-16'h015c,16'h020f,16'h000b,16'h0070,-16'h019c,16'h01da,-16'h002b,-16'h0182,-16'h016c,-16'h00e1,16'h0046,16'h014a,-16'h0387,16'h0044,-16'h0062,-16'h0090,16'h00e9,16'h00ff,-16'h004a,16'h0012,16'h00fa,16'h0071,16'h00a8,-16'h0079,16'h001d,-16'h0380,-16'h0124,-16'h005e,-16'h0061,16'h00ce,-16'h016b,-16'h0456,-16'h00bf,-16'h003e,-16'h00b5,16'h003d,16'h0169,-16'h0032,-16'h00d5,16'h00e7,16'h00ce,-16'h003b,-16'h00d6,-16'h00b4,16'h018b,16'h0099,-16'h006e,-16'h0026,-16'h013e,-16'h002c,16'h0066,16'h003f,16'h013d,-16'h0139,16'h0039,-16'h014b,16'h0002,16'h007b,-16'h0176,16'h0112,16'h0045,16'h0007,-16'h006f,-16'h0003,-16'h022c,16'h023d,16'h000e,-16'h0012,-16'h00ec,16'h01a7,-16'h0011,16'h0000,-16'h0173,-16'h00bb,16'h0007,16'h006a,-16'h03ee,16'h0122,-16'h00c1,-16'h0145,16'h0144,16'h0114,-16'h003a,16'h008f,16'h0078,16'h0069,16'h0031,-16'h00e1,16'h0026,-16'h0544,-16'h0122,-16'h00a8,16'h0043,16'h00c6,-16'h00ff,-16'h0362,-16'h0103,16'h0080,-16'h00b5,16'h0027,16'h0113,-16'h02a9,-16'h0098,16'h0091,16'h006e,-16'h0121,-16'h0078,-16'h0113,16'h00b4,16'h00a6,-16'h0316,16'h005b,-16'h0008,-16'h0012,16'h0102,16'h0078,16'h0172,-16'h0047,16'h007b,-16'h0100,16'h0062,16'h008f,-16'h012b,16'h0085,16'h0102,16'h0015,-16'h0025,-16'h0040,-16'h023f,16'h01b6,16'h0080,-16'h0075,-16'h00aa,16'h0010,16'h006b,16'h00e4,-16'h0161,-16'h0107,16'h007d,-16'h0070,-16'h0340,16'h0140,-16'h00d4,-16'h00b6,16'h01a0,16'h0184,-16'h0039,16'h008c,16'h0092,-16'h003e,16'h0040,-16'h0051,16'h002d,-16'h054f,-16'h0169,-16'h00a4,-16'h0020,16'h0150,-16'h00fa,-16'h026b,-16'h00f2,16'h00b0,-16'h00a9,16'h0037,16'h0106,-16'h04ea,-16'h003f,16'h0082,-16'h004f,-16'h0280,-16'h000c,-16'h010a,-16'h003b,16'h004e,-16'h0274,16'h0009,16'h01e1,-16'h0068,16'h007b,16'h0060,16'h0148,16'h002a,-16'h00bd,-16'h0139,16'h006f,16'h0000,-16'h00d6,-16'h0018,16'h0041,16'h0034,-16'h0035,-16'h00ae,-16'h0168,16'h0121,-16'h0015,16'h003f,-16'h00eb,-16'h01ce,16'h0050,16'h00c1,-16'h00e9,-16'h00a7,16'h0006,-16'h0088,-16'h031a,16'h0144,-16'h0043,-16'h00bb,16'h0115,16'h0170,-16'h007b,16'h00d5,16'h007b,-16'h0020,16'h004c,16'h0008,16'h0010,-16'h0394,-16'h006f,16'h0027,-16'h0003,16'h00fb,16'h0006,-16'h01d0,-16'h012c,16'h000a,-16'h009a,-16'h0026,16'h00fc,-16'h0511,-16'h00b2,-16'h0086,-16'h01b9,-16'h029f,-16'h000f,-16'h0179,-16'h0228,16'h007f,-16'h00a2,-16'h0047,16'h02d7,16'h0057,16'h0015,16'h0048,16'h017b,-16'h0061,-16'h0165,-16'h0116,16'h0077,16'h00ae,-16'h0101,-16'h0060,16'h014c,-16'h0015,-16'h0022,-16'h007b,-16'h009c,16'h006e,16'h0026,16'h0099,-16'h014e,-16'h0198,16'h009c,16'h004c,-16'h00cc,16'h0030,-16'h001e,-16'h0158,-16'h0301,16'h00db,-16'h00a2,16'h0006,16'h0039,16'h0169,-16'h0029,16'h009c,16'h0083,-16'h002e,16'h0119,16'h0071,16'h001d,-16'h00a3,16'h0009,16'h0145,16'h0010,16'h00f5,-16'h0041,-16'h00c6,-16'h0065,-16'h000f,-16'h007a,16'h006c,16'h0139,-16'h037f,-16'h005b,-16'h0132,-16'h048b,-16'h019b,16'h007e,-16'h0239,-16'h02d9,-16'h0058,16'h00fa,16'h00bc,16'h01c1,16'h0011,-16'h0059,16'h008c,16'h019b,16'h0070,-16'h00fc,-16'h0115,16'h006e,16'h0138,-16'h010d,16'h000f,16'h01a0,-16'h0074,16'h0059,-16'h0101,-16'h0041,16'h007b,16'h0037,16'h00fb,-16'h00a9,-16'h0202,-16'h0003,-16'h0010,-16'h00c5,16'h0092,16'h0152,-16'h012a,-16'h035d,16'h00fa,-16'h005d,-16'h0119,16'h006d,16'h0129,16'h0053,16'h0056,16'h00a1,-16'h002d,16'h0083,16'h0078,-16'h0042,16'h0170,-16'h0122,16'h0256,-16'h0117,16'h000e,16'h007d,-16'h006d,-16'h00b7,-16'h011e,16'h0019,16'h0105,16'h01ad,-16'h01ef,-16'h00d9,-16'h011f,-16'h04b9,-16'h002b,-16'h0011,-16'h02ba,-16'h0378,-16'h0099,16'h014b,16'h0155,16'h002c,-16'h0081,-16'h0107,16'h0196,16'h0158,16'h0162,-16'h0065,-16'h00ab,16'h00d0,16'h018d,-16'h0113,16'h009a,16'h011a,-16'h0002,-16'h0089,-16'h001f,-16'h00de,16'h0083,16'h0003,16'h0185,-16'h00bb,-16'h014a,-16'h00b9,-16'h00c2,-16'h0056,16'h001c,16'h01e7,-16'h01b8,-16'h0347,16'h00d0,-16'h0114,-16'h0292,16'h00a5,16'h016d,16'h0042,16'h0128,16'h0088,-16'h00fc,16'h0132,-16'h002f,-16'h000f,16'h029d,-16'h022a,16'h014b,-16'h01c1,-16'h0092,16'h012f,-16'h000f,-16'h01e5,-16'h0177,-16'h0039,16'h00e8,16'h018f,-16'h0068,-16'h01f3,-16'h005b,-16'h0380,16'h0037,16'h000d,-16'h032b,-16'h01c8,-16'h002c,16'h0128,16'h0232,16'h002e,-16'h011c,-16'h01b3,16'h021b,16'h0273,16'h01bd,-16'h00f7,-16'h016d,16'h00d0,16'h01a5,-16'h0054,-16'h0006,-16'h005c,-16'h00e8,-16'h00e0,-16'h002f,-16'h013d,16'h001e,-16'h0015,16'h026f,-16'h00f7,-16'h0071,16'h0004,-16'h01fd,-16'h00d6,-16'h008b,16'h0185,-16'h007d,-16'h0001,-16'h0199,-16'h0127,-16'h00df,-16'h00b3,16'h0125,-16'h00f0,16'h001b,-16'h009c,16'h00ae,16'h0336,-16'h008f,16'h008c,16'h0101,16'h00c3,16'h0012,-16'h0051,-16'h00b0,-16'h0018,16'h002a,16'h0021,16'h004b,16'h0057,-16'h0070,-16'h00ac,16'h004e,16'h0089,-16'h0049,16'h0065,16'h0046,-16'h0010,16'h010a,-16'h00bf,16'h008e,-16'h0009,-16'h009b,-16'h0036,-16'h00aa,16'h01dd,-16'h00e4,16'h002e,16'h015e,16'h0166,16'h002b,-16'h00b0,16'h0009,-16'h015c,16'h0019,16'h00b3,-16'h003c,-16'h0045,-16'h0052,-16'h01a3,-16'h00a1,16'h0145,16'h010a,16'h00c8,-16'h0014,-16'h00b9,16'h0098,16'h00e1,16'h0034,16'h01bd,-16'h005d,16'h0020,-16'h0146,-16'h019f,-16'h0082,16'h0004,16'h0198,-16'h013d,16'h0086,-16'h0083,-16'h0084,16'h02b8,-16'h0070,16'h015a,16'h000e,16'h0152,16'h003e,-16'h002c,-16'h000b,16'h003b,16'h006a,-16'h00da,-16'h00d3,-16'h0043,16'h0029,-16'h0031,-16'h0040,-16'h0047,-16'h0093,16'h004c,16'h00ff,16'h006e,16'h00ff,-16'h0066,-16'h0032,16'h005b,-16'h0044,16'h0012,-16'h0027,16'h0183,-16'h0073,16'h004e,16'h013a,16'h00ec,-16'h0038,-16'h0009,16'h0093,-16'h00ea,-16'h0009,16'h00e5,-16'h008c,16'h0054,-16'h0007,16'h000d,-16'h0069,16'h0111,16'h00cd,16'h0107,16'h00ab,-16'h008c,16'h0149,16'h00ed,16'h0014,16'h01cd,-16'h0042,16'h0022,-16'h00f1,-16'h020a,-16'h0059,16'h0079,16'h015e,-16'h0098,16'h0093,-16'h00ad,-16'h0163,16'h01b9,-16'h0048,16'h015d,16'h000f,16'h0138,16'h0066,-16'h00e6,16'h009f,16'h006c,16'h0089,-16'h01f0,-16'h0143,-16'h0006,16'h00b1,-16'h0062,16'h0039,-16'h0038,-16'h0092,16'h0076,16'h006c,16'h00d5,16'h0061,16'h0070,-16'h00a5,16'h000d,-16'h0113,16'h0006,-16'h012d,16'h0194,-16'h0094,-16'h001b,16'h0170,16'h00fe,-16'h0035,16'h001f,-16'h002a,-16'h0008,-16'h0048,16'h00c8,-16'h012d,16'h005a,16'h0021,16'h000f,-16'h00bf,16'h00fd,16'h013a,16'h0053,16'h009f,-16'h0094,16'h0105,16'h0116,-16'h0027,16'h00e1,-16'h0037,16'h0045,16'h0002,-16'h0299,-16'h006d,16'h00bf,16'h00ca,-16'h0038,16'h00a9,-16'h0042,-16'h01aa,16'h01e3,-16'h003e,16'h002e,-16'h0020,16'h01b5,16'h0089,-16'h0040,16'h013f,16'h011f,16'h0130,-16'h01f8,-16'h014a,-16'h004d,16'h0062,-16'h00dc,-16'h000b,-16'h006e,-16'h0035,-16'h0054,16'h00cd,16'h002a,16'h0011,16'h00a1,-16'h00d7,16'h006b,-16'h0082,-16'h0068,-16'h0146,16'h01b2,-16'h0039,16'h0070,16'h0061,16'h015e,16'h001e,16'h0063,16'h0069,16'h0083,16'h0023,16'h00d6,-16'h0116,-16'h0073,16'h0039,16'h0027,-16'h0182,16'h012c,16'h00a0,16'h0076,16'h0062,-16'h003f,16'h00e1,16'h011c,-16'h0082,16'h00fa,-16'h0029,-16'h0047,16'h002b,-16'h031c,-16'h0027,-16'h0007,16'h00c5,16'h0013,16'h0049,-16'h0041,-16'h01b0,16'h0145,-16'h0052,-16'h0056,16'h0004,16'h00e7,16'h0071,-16'h0010,16'h0180,16'h0119,16'h00b3,-16'h0265,-16'h0201,16'h003f,16'h006f,16'h0074,-16'h0031,-16'h0064,16'h0038,-16'h0089,16'h0103,16'h00a9,16'h0002,16'h0100,-16'h00f3,16'h0030,-16'h00a0,-16'h00f9,-16'h01a5,16'h013b,-16'h0046,16'h00cd,-16'h0102,16'h00f8,16'h00cf,16'h00ad,16'h00b9,16'h00bb,16'h00b4,16'h0137,-16'h0088,-16'h003a,-16'h0051,-16'h0012,-16'h01a1,16'h0036,16'h0120,16'h00ea,16'h0023,16'h0028,16'h006f,16'h0136,-16'h0089,16'h0090,16'h0060,16'h0059,16'h008b,-16'h0333,-16'h00a1,16'h008d,16'h0098,16'h0051,16'h0025,-16'h005e,-16'h0145,16'h014a,16'h0030,-16'h01bf,16'h0082,16'h00e7,16'h001c,-16'h0022,16'h0168,16'h0080,16'h00ad,-16'h019c,-16'h0128,16'h0000,-16'h00fb,16'h00a6,-16'h000c,-16'h0071,16'h0061,-16'h00a4,16'h00c2,16'h006a,-16'h008e,16'h006a,16'h0000,16'h007a,-16'h009b,16'h001a,-16'h00fc,16'h00f3,-16'h006e,16'h00bf,-16'h0155,16'h0091,16'h00d0,-16'h003a,16'h0038,16'h004c,16'h00eb,16'h011a,-16'h0090,16'h001d,-16'h0038,-16'h0004,-16'h0229,-16'h0028,16'h0093,16'h0066,16'h00bb,16'h005f,16'h00f2,16'h00f0,16'h00be,16'h0105,16'h00a8,16'h002b,-16'h0041,-16'h02c9,-16'h00de,-16'h0012,16'h00e0,16'h002e,-16'h005a,-16'h0078,-16'h00d3,16'h0057,16'h0056,-16'h018d,16'h00be,16'h00ba,-16'h001e,16'h0081,16'h021e,16'h001f,16'h0045,-16'h015a,16'h0032,-16'h0007,-16'h00d1,16'h00ab,-16'h008d,-16'h00c5,16'h00ec,-16'h0060,16'h00fe,-16'h00fa,-16'h00f9,-16'h0053,16'h0126,16'h00a9,-16'h00bb,-16'h001b,-16'h010b,16'h014b,-16'h007b,16'h016a,-16'h0223,-16'h0005,16'h00a2,-16'h008b,16'h00bc,-16'h001d,16'h00ee,16'h00eb,-16'h00bc,16'h0008,16'h000e,16'h004e,-16'h0160,-16'h0103,16'h0099,16'h0070,16'h00f7,16'h000a,16'h0093,16'h00de,16'h0154,16'h00ba,16'h001f,-16'h002b,-16'h0044,-16'h0284,-16'h0107,16'h00b1,16'h00f4,16'h003c,-16'h001e,-16'h00c7,-16'h01b5,-16'h0036,16'h003d,16'h0072,16'h00bf,16'h00c2,16'h004d,16'h0024,16'h0179,-16'h003d,-16'h007d,-16'h00fb,16'h00f6,-16'h006b,-16'h00c9,-16'h0028,-16'h010f,-16'h00a2,-16'h0013,-16'h003a,16'h00c0,-16'h01f9,-16'h00b5,16'h0021,16'h0138,-16'h000c,-16'h0067,16'h0058,-16'h00a7,16'h003d,-16'h007f,16'h01b4,-16'h023e,16'h008a,-16'h0002,-16'h00c6,16'h00da,-16'h00b4,16'h0023,16'h0139,-16'h00e3,16'h00b0,-16'h0064,16'h0052,-16'h01e6,-16'h01db,-16'h0018,16'h00ba,16'h00f2,-16'h008a,16'h0094,16'h00fd,16'h010a,16'h008e,16'h000c,-16'h0093,-16'h017c,-16'h01ce,-16'h00d4,16'h003f,16'h00c0,16'h0063,16'h0022,-16'h005e,-16'h01c8,-16'h003b,-16'h008f,16'h023e,16'h0166,16'h0064,16'h0108,16'h0004,16'h018d,16'h001e,-16'h00d8,-16'h000e,16'h00af,-16'h00f8,-16'h008e,-16'h0047,-16'h0123,-16'h0093,-16'h0022,-16'h0049,16'h00e9,-16'h032c,-16'h0198,-16'h0002,-16'h0020,-16'h006c,-16'h0080,-16'h0068,-16'h0131,16'h0043,-16'h00d2,16'h0121,-16'h01c2,16'h0109,16'h001a,-16'h002e,16'h01b7,-16'h00c0,-16'h00a6,16'h00d9,-16'h0053,16'h00bb,-16'h0126,-16'h0018,-16'h01bb,-16'h0184,16'h002d,16'h0059,16'h00ad,16'h0041,16'h0032,16'h0106,16'h017e,16'h006b,-16'h002c,-16'h012b,-16'h0178,-16'h0222,-16'h00cc,16'h0078,16'h0129,16'h0038,16'h0078,-16'h014b,-16'h0241,-16'h012e,-16'h0010,16'h0230,16'h0138,16'h0040,16'h00fb,16'h0099,16'h01bb,16'h0070,-16'h0193,16'h0103,16'h0096,-16'h00ea,16'h0158,-16'h00cd,-16'h00e0,-16'h00bd,-16'h005a,16'h003d,16'h007a,-16'h031e,-16'h01a1,16'h00dc,-16'h01ba,-16'h0061,-16'h0030,16'h00a7,-16'h011f,-16'h0001,16'h0013,16'h0091,-16'h012e,16'h0101,-16'h001d,16'h006f,16'h0133,-16'h0121,-16'h0086,16'h0192,16'h008c,16'h0089,-16'h00d5,-16'h0027,-16'h0189,16'h007f,-16'h0032,-16'h0088,16'h0111,16'h00b8,16'h003d,16'h00a2,16'h01b8,-16'h00eb,-16'h0080,-16'h011f,-16'h00f0,-16'h0140,-16'h0015,16'h0078,16'h00d7,16'h0069,16'h00c1,-16'h00d0,-16'h025e,-16'h026a,-16'h000e,16'h0152,16'h0085,16'h0045,16'h0111,-16'h002a,16'h01ea,16'h00c7,-16'h00d3,16'h018c,16'h0085,-16'h0167,16'h0208,-16'h006f,-16'h00cf,-16'h0078,-16'h0064,16'h0037,16'h0166,-16'h0193,-16'h016c,16'h013e,-16'h0307,16'h0110,-16'h006a,16'h007a,-16'h0129,16'h0082,16'h0061,16'h00ad,-16'h00ae,16'h00bd,16'h0026,16'h0067,16'h0138,-16'h0136,-16'h0055,16'h015c,16'h0034,16'h00f5,-16'h006b,-16'h0049,-16'h00d1,16'h0111,-16'h0004,16'h0004,16'h018c,-16'h0010,16'h0036,16'h00df,16'h00c5,-16'h0042,-16'h007d,-16'h0097,-16'h00ec,-16'h014a,-16'h0043,16'h00b3,16'h00e0,16'h0107,16'h0059,-16'h003e,-16'h0245,-16'h01b8,16'h0022,-16'h00ff,-16'h00d9,16'h0047,16'h00a5,16'h0014,16'h01da,16'h0126,16'h0039,16'h010b,16'h006c,-16'h0169,16'h02b7,-16'h00b5,-16'h00b2,-16'h00ae,16'h006a,-16'h008c,16'h011d,16'h0037,-16'h0248,16'h00e0,-16'h02ba,16'h0221,16'h0013,-16'h006c,-16'h0120,16'h00ce,-16'h0009,-16'h002e,16'h003e,16'h00cc,16'h0077,16'h0099,16'h0080,-16'h01b0,-16'h0028,16'h0191,16'h000c,16'h0111,16'h005f,16'h007f,-16'h00f8,16'h00da,16'h006e,-16'h002c,16'h0125,-16'h0034,16'h006e,16'h0086,16'h015a,-16'h0041,16'h001e,-16'h0092,-16'h015b,-16'h0112,-16'h00b9,16'h00e3,16'h0192,16'h0026,16'h0111,-16'h0045,-16'h01b6,-16'h01cc,16'h0047,-16'h0154,-16'h0111,-16'h003a,16'h0031,-16'h0089,16'h0277,16'h010a,16'h0096,16'h00bc,-16'h002a,-16'h00fa,16'h01e2,-16'h00df,-16'h009c,-16'h00c0,16'h00eb,-16'h012b,-16'h0075,16'h00c4,-16'h01bc,16'h0110,-16'h004f,16'h0220,16'h0013,-16'h0172,-16'h00fb,16'h0164,-16'h0003,-16'h007e,16'h00ab,16'h0050,16'h0062,16'h00e6,16'h007c,-16'h01c7,-16'h0016,16'h014f,16'h00fc,16'h00e8,16'h003d,16'h0122,-16'h008e,16'h011f,16'h0037,-16'h0010,16'h0091,-16'h002d,16'h002a,16'h008a,16'h016a,-16'h0067,16'h00ba,-16'h00a2,-16'h0186,-16'h010e,-16'h018c,16'h00e7,16'h0156,-16'h00e7,16'h0029,-16'h0008,-16'h018f,-16'h00f2,16'h002c,-16'h011c,-16'h0105,-16'h001c,16'h0081,-16'h00bf,16'h0264,16'h0091,16'h006c,16'h00d4,-16'h00cf,-16'h00c5,16'h01f4,-16'h0094,16'h000f,-16'h00bd,16'h01e4,-16'h0133,-16'h00b9,16'h013d,-16'h0132,16'h0141,16'h007d,-16'h0089,-16'h0081,16'h002d,-16'h0124,16'h00d7,-16'h0089,-16'h0012,16'h00d2,16'h005e,-16'h0066,16'h0078,-16'h0001,-16'h0251,16'h0029,16'h0189,16'h0137,16'h004d,16'h0040,16'h00f1,-16'h0071,16'h00bd,16'h00d9,16'h0002,16'h008c,-16'h001e,-16'h0008,16'h0007,16'h01ef,-16'h003a,16'h0007,-16'h004e,-16'h0131,-16'h0129,-16'h0247,16'h01a4,16'h0114,-16'h013e,-16'h0032,-16'h00af,-16'h0160,16'h008a,16'h000a,16'h0085,-16'h008d,-16'h0060,16'h0073,-16'h00ab,16'h0218,16'h0084,16'h0074,16'h0099,-16'h00af,-16'h00ea,16'h00ca,-16'h007a,16'h005a,-16'h00c0,16'h0195,-16'h008e,-16'h0045,16'h0132,-16'h0130,-16'h0045,16'h0016,-16'h0295,16'h0001,16'h00f8,-16'h019a,16'h00be,-16'h0041,-16'h005d,16'h00c2,16'h0065,-16'h008a,16'h00e2,16'h002b,-16'h0213,-16'h001d,16'h01ce,16'h005d,16'h009d,16'h00ac,16'h00d6,16'h0007,-16'h000b,16'h006b,16'h0029,16'h009b,-16'h007d,-16'h0086,-16'h006e,16'h0203,-16'h0027,16'h0080,-16'h006a,-16'h0092,-16'h011f,-16'h0222,16'h0179,16'h00d0,-16'h0091,-16'h00aa,-16'h00ef,-16'h0009,16'h010c,16'h004e,16'h014e,16'h0023,-16'h0052,16'h009e,-16'h00e7,16'h0186,16'h0087,-16'h000f,16'h006f,-16'h00ee,-16'h00af,-16'h00e2,-16'h003c,-16'h0019,-16'h00c9,16'h0168,-16'h00a8,-16'h006c,16'h015f,-16'h012d,-16'h01f9,16'h008f,-16'h01f4,16'h0052,16'h002b,-16'h00e9,16'h0004,-16'h009d,-16'h0110,16'h001b,16'h0065,-16'h0030,16'h023d,16'h0007,-16'h016c,-16'h00a5,16'h018b,16'h000a,16'h0029,16'h0043,16'h015f,16'h0095,16'h004f,16'h004d,16'h0047,16'h00ab,-16'h0093,-16'h0108,-16'h0020,16'h01a9,-16'h0036,16'h00c0,-16'h015c,-16'h013d,-16'h00e4,-16'h0224,16'h024f,16'h0105,-16'h019b,16'h0004,-16'h00b4,16'h00a8,16'h00cb,16'h0000,16'h0114,16'h0032,-16'h00df,16'h00a0,-16'h00cd,16'h0174,16'h00da,16'h0033,16'h00b9,-16'h012b,-16'h00f2,-16'h014b,-16'h000f,16'h003f,-16'h0110,16'h0052,-16'h000a,-16'h0041,16'h014b,-16'h00d7,-16'h0322,16'h00be,-16'h005f,16'h0083,-16'h0023,-16'h0078,-16'h0059,-16'h0024,-16'h0090,-16'h008a,16'h0009,16'h0009,16'h01c1,16'h005e,-16'h0159,-16'h0114,16'h0155,-16'h0025,16'h0012,16'h0016,16'h008e,16'h00ff,-16'h004c,16'h00a3,-16'h0014,16'h0069,-16'h000f,-16'h016e,-16'h0025,16'h0088,16'h002a,16'h00bd,-16'h01d3,-16'h007f,-16'h011c,-16'h01ee,16'h0215,16'h00d7,-16'h0161,16'h00cc,16'h005a,16'h0066,16'h003c,16'h005f,16'h00d3,16'h002f,16'h0024,16'h007c,-16'h012b,16'h017c,16'h00b7,16'h000c,16'h0085,-16'h00b6,-16'h013a,-16'h002f,-16'h0013,16'h0057,-16'h0084,-16'h0003,16'h007c,16'h008e,16'h0052,-16'h010d,-16'h02d4,16'h005d,16'h00a0,16'h004c,-16'h0005,-16'h001b,-16'h0145,-16'h004c,-16'h0010,-16'h00c3,-16'h0071,16'h0039,16'h00d8,16'h0093,-16'h0155,-16'h00b4,16'h018e,16'h005c,16'h0008,16'h007e,-16'h002c,16'h0147,-16'h0029,16'h0008,-16'h0042,16'h012c,16'h0005,-16'h0191,-16'h00ba,16'h009a,16'h0042,16'h0113,-16'h016b,-16'h0037,-16'h0186,-16'h0145,16'h019d,16'h00f4,-16'h00f7,16'h00e3,16'h009b,16'h003c,16'h0009,-16'h0048,16'h008d,16'h0121,-16'h0006,16'h011d,-16'h0051,16'h00f3,16'h00b8,-16'h00b4,-16'h0088,-16'h0090,-16'h00e0,-16'h00c4,16'h0040,16'h004d,-16'h00f6,-16'h0097,16'h00d1,16'h0089,16'h003b,-16'h00d5,-16'h010d,16'h0096,16'h0132,-16'h0017,-16'h0052,-16'h000e,-16'h010f,-16'h0048,16'h0062,-16'h0081,16'h0047,-16'h00f9,16'h005c,16'h0046,-16'h014c,-16'h0040,16'h017b,16'h00b0,-16'h0002,16'h003e,-16'h013d,16'h0116,-16'h0072,16'h00c0,-16'h005b,16'h00af,-16'h0031,-16'h02a8,-16'h00a3,-16'h0022,16'h0095,16'h014e,-16'h024b,-16'h00b1,-16'h00ff,-16'h00ea,16'h019e,16'h0135,-16'h0088,16'h017e,16'h00d0,16'h002b,16'h000c,16'h0012,16'h0066,16'h010f,16'h000b,16'h009f,-16'h00a8,16'h0141,-16'h0054,-16'h0173,-16'h001f,-16'h0016,-16'h0142,-16'h00e8,16'h00c5,-16'h0075,-16'h012c,16'h008d,16'h008d,16'h00a3,16'h0015,-16'h00cc,16'h003b,16'h0029,16'h00e9,-16'h0032,-16'h00fc,-16'h0008,16'h001f,-16'h0028,16'h009a,-16'h011e,16'h002b,-16'h0136,-16'h001d,-16'h0007,-16'h00bf,16'h0091,16'h00d8,16'h008c,-16'h0063,16'h0035,-16'h015d,16'h0146,-16'h0044,16'h00e9,-16'h0100,16'h0158,-16'h001f,-16'h029d,-16'h0057,-16'h012b,16'h0041,16'h0111,-16'h0323,-16'h004f,-16'h013a,-16'h00e3,16'h0130,16'h0098,-16'h00ef,16'h0063,16'h0140,16'h00a2,16'h00a3,-16'h0053,16'h001f,-16'h006d,-16'h00cd,16'h00b1,-16'h0077,16'h00d6,-16'h0099,-16'h03fe,-16'h00b4,-16'h0090,-16'h0065,-16'h0098,16'h0115,-16'h004d,-16'h00d0,16'h00ff,16'h0140,16'h002c,-16'h0047,-16'h00aa,16'h01b9,16'h001d,16'h0032,-16'h0035,-16'h0158,16'h0039,-16'h000e,16'h0063,16'h00e7,-16'h01a6,16'h00c1,-16'h00cd,-16'h0015,16'h0052,-16'h013f,16'h00be,-16'h002d,16'h0065,-16'h003f,-16'h0023,-16'h0160,16'h0153,16'h0079,16'h009e,-16'h0092,16'h0121,-16'h0082,-16'h0261,-16'h014e,-16'h0255,-16'h0063,16'h018e,-16'h0443,-16'h0062,-16'h018b,-16'h00c1,16'h018a,16'h00b8,-16'h0147,16'h003e,16'h012f,16'h0095,16'h0122,-16'h00a6,-16'h0008,-16'h02f4,-16'h00f0,16'h006d,-16'h0066,16'h0096,-16'h0143,-16'h04fd,-16'h0166,-16'h0060,-16'h00ab,16'h00b9,16'h0178,-16'h017d,-16'h0071,16'h011a,16'h00d9,-16'h0110,-16'h0057,-16'h00ad,16'h0186,-16'h0034,-16'h017a,-16'h0058,-16'h0068,16'h006f,16'h002b,16'h005a,16'h0199,-16'h014c,16'h0136,-16'h00dd,-16'h0041,16'h0031,-16'h0208,16'h0097,16'h006f,16'h0088,16'h0001,-16'h0049,-16'h01bc,16'h0199,16'h0092,16'h0050,-16'h0006,-16'h0049,16'h0055,-16'h009d,-16'h0150,-16'h0301,-16'h003b,16'h00fa,-16'h040b,16'h0075,-16'h01bf,-16'h011f,16'h017b,16'h0137,-16'h00b4,16'h0061,16'h0112,16'h0087,16'h010f,-16'h0036,-16'h0048,-16'h0517,-16'h01e0,16'h0041,16'h0037,16'h0076,-16'h010a,-16'h03e2,-16'h01a1,16'h008b,-16'h0097,16'h004f,16'h011a,-16'h03d5,-16'h00dd,16'h00a6,16'h0046,-16'h0185,16'h0028,-16'h00d3,16'h00c2,-16'h0088,-16'h02d7,-16'h0067,16'h005e,16'h009d,16'h00c2,16'h00ab,16'h013f,-16'h0044,16'h00e6,-16'h009f,16'h00ab,16'h0046,-16'h01d6,16'h00bf,16'h0077,16'h001d,-16'h004b,-16'h003d,-16'h01c2,16'h0188,16'h00b5,16'h0009,-16'h00b2,-16'h011a,16'h0036,16'h00de,-16'h00a1,-16'h01e7,16'h004b,16'h007e,-16'h02d4,16'h004c,-16'h0234,-16'h00c3,16'h013e,16'h016f,-16'h00b8,16'h007f,16'h00ee,16'h0058,16'h006e,-16'h0040,-16'h0029,-16'h04b8,-16'h015b,-16'h000e,-16'h000a,16'h00cf,-16'h009d,-16'h0306,-16'h0169,16'h006c,-16'h00c3,16'h0072,16'h0103,-16'h0519,-16'h00fa,16'h000e,-16'h000d,-16'h034c,16'h005b,-16'h00b5,-16'h00d4,-16'h0046,-16'h0297,-16'h00ac,16'h026f,16'h0093,16'h0067,16'h0087,16'h016f,16'h0078,16'h0035,-16'h00a5,16'h00d3,16'h00e8,-16'h0164,-16'h0025,16'h0082,-16'h0031,16'h0018,-16'h002e,-16'h0133,16'h00be,16'h0045,16'h003f,-16'h004f,-16'h01d2,-16'h000e,16'h00ff,-16'h00da,-16'h006a,-16'h0007,16'h0059,-16'h0279,16'h00e6,-16'h01c5,-16'h00c8,16'h00f6,16'h017e,-16'h0027,16'h005d,16'h00a2,-16'h001e,16'h0076,-16'h000d,16'h0075,-16'h03b6,-16'h003f,-16'h000d,16'h0055,16'h00fe,-16'h0066,-16'h0211,-16'h0214,16'h004a,-16'h0110,16'h0011,16'h015c,-16'h041d,-16'h00da,-16'h0096,-16'h023f,-16'h03df,16'h0068,-16'h0128,-16'h0332,16'h0053,-16'h006c,16'h0019,16'h025c,16'h0035,-16'h0042,16'h0062,16'h00d1,-16'h0016,-16'h00ba,-16'h00a3,16'h00cc,16'h00c5,-16'h00f6,-16'h002d,16'h00ef,-16'h0033,16'h0041,16'h008e,-16'h0050,16'h003b,16'h0014,16'h004c,-16'h0063,-16'h0120,16'h002a,16'h0121,-16'h00fe,-16'h0004,16'h000c,-16'h009c,-16'h02ba,16'h00a5,-16'h00ac,16'h0016,16'h006d,16'h00d1,16'h0090,16'h0010,16'h007e,16'h0000,16'h00cb,16'h008d,-16'h0093,-16'h00dc,16'h0029,16'h0135,16'h008b,16'h00ac,-16'h002d,-16'h0137,-16'h00c8,-16'h0035,-16'h017a,16'h00b7,16'h0204,-16'h037a,-16'h005b,-16'h0136,-16'h0587,-16'h0246,16'h00a2,-16'h021a,-16'h03e8,-16'h008f,16'h00e1,16'h00ad,16'h0169,16'h0002,-16'h0011,16'h009f,16'h0141,16'h0067,-16'h0089,-16'h001f,16'h003f,16'h014b,-16'h00f3,-16'h001c,16'h0172,-16'h0070,16'h0021,16'h0003,-16'h005e,16'h0063,-16'h0032,16'h00df,-16'h009e,-16'h0177,-16'h0056,16'h0024,-16'h006e,16'h0048,16'h017f,-16'h012f,-16'h035f,16'h0080,-16'h00f1,-16'h005b,16'h00af,16'h010e,16'h00ba,-16'h004f,16'h00ef,-16'h002d,-16'h0049,16'h005c,-16'h006f,16'h01b1,-16'h0126,16'h024a,-16'h0122,16'h0099,-16'h0036,-16'h004f,-16'h010a,-16'h00bc,-16'h013b,16'h0103,16'h01a4,-16'h01cf,-16'h00b8,-16'h015f,-16'h04b0,-16'h011c,16'h00b1,-16'h02f8,-16'h038c,-16'h0084,16'h0159,16'h0102,16'h004e,-16'h004d,-16'h0026,16'h0169,16'h00e2,16'h011a,-16'h00b1,-16'h0043,16'h0163,16'h00f8,-16'h006f,-16'h001f,16'h00f6,16'h0018,16'h0010,16'h005e,-16'h0054,-16'h003c,16'h006d,16'h00d8,-16'h004e,-16'h0086,-16'h0161,-16'h0144,-16'h0045,16'h0048,16'h0250,-16'h0169,-16'h0360,16'h0080,-16'h0102,-16'h01a2,16'h0066,16'h00ad,16'h003d,16'h0002,16'h00cd,-16'h011c,16'h0118,-16'h004a,-16'h0018,16'h0285,-16'h0279,16'h0145,-16'h0269,-16'h000a,16'h0082,-16'h0065,-16'h0147,-16'h0190,-16'h0179,16'h0122,16'h01c1,16'h0030,-16'h023e,-16'h005a,-16'h03e9,-16'h004d,16'h0030,-16'h0320,-16'h023c,16'h007a,16'h01e4,16'h0195,-16'h00aa,-16'h01a0,-16'h0109,16'h0268,16'h011a,16'h0156,-16'h0087,-16'h00c6,16'h01bb,16'h0149,-16'h002a,-16'h002f,-16'h0075,-16'h0024,-16'h0127,16'h0016,-16'h0147,-16'h010e,16'h0028,16'h0278,-16'h00d2,-16'h00a5,-16'h00b1,-16'h02d1,-16'h005e,-16'h012b,16'h015b,-16'h0068,16'h00bb,-16'h01c6,-16'h010b,-16'h0079,-16'h0075,16'h00a1,-16'h0031,-16'h0025,-16'h012c,16'h0096,16'h02f9,-16'h004a,16'h00b8,16'h00a5,16'h00db,-16'h0113,-16'h0004,-16'h0118,16'h006a,-16'h007e,-16'h0097,-16'h0023,16'h0054,-16'h00a1,-16'h0183,-16'h00be,16'h00bb,-16'h00a2,16'h0117,16'h00cd,16'h004c,16'h0163,16'h0020,16'h00bb,-16'h0048,16'h0058,16'h0092,-16'h0145,16'h01ad,-16'h009c,16'h002f,16'h00b8,16'h01a5,16'h00a0,-16'h0111,16'h0089,-16'h0160,16'h0015,16'h00b2,-16'h001d,-16'h0088,-16'h0067,-16'h01ae,-16'h01d5,16'h017c,16'h00a9,16'h00ff,16'h004e,-16'h006a,16'h00d8,-16'h0018,-16'h00e7,16'h01c8,-16'h007b,16'h0038,-16'h012c,-16'h015a,-16'h0013,16'h002d,16'h0118,-16'h009b,16'h0038,-16'h00d2,-16'h0067,16'h02a0,-16'h00e7,16'h00f0,16'h000c,16'h00b0,-16'h00ba,-16'h002a,-16'h00e3,16'h00a8,-16'h009c,-16'h00ae,-16'h014e,16'h0052,16'h0043,-16'h00dd,-16'h00c4,16'h000c,-16'h0027,16'h0068,16'h00d4,16'h0049,16'h013f,16'h001a,16'h0018,16'h0014,16'h0034,-16'h0067,-16'h015e,16'h01bf,-16'h0092,16'h0067,16'h015e,16'h0133,-16'h004a,-16'h001c,16'h0083,-16'h00ae,-16'h004d,16'h00a9,-16'h011b,-16'h0006,-16'h0036,-16'h011a,-16'h0186,16'h0112,16'h00be,16'h00a4,16'h0009,-16'h006e,16'h0126,16'h0079,-16'h0091,16'h011b,16'h004d,16'h0006,-16'h014c,-16'h024f,16'h0022,16'h005c,16'h0094,-16'h00e9,16'h005d,-16'h0132,-16'h0139,16'h023b,-16'h006a,16'h011f,-16'h004c,16'h0123,-16'h00df,16'h000c,-16'h0071,16'h005b,16'h0063,-16'h0184,-16'h00a2,-16'h0017,16'h0050,-16'h0125,-16'h00a8,-16'h0013,-16'h000d,16'h001f,16'h0100,16'h00d6,16'h0127,16'h0084,-16'h0089,16'h0000,-16'h005d,-16'h0005,-16'h01e1,16'h020b,-16'h004a,-16'h0011,16'h010d,16'h00a8,16'h0073,16'h001e,16'h0080,-16'h0070,16'h0032,16'h006c,-16'h008c,16'h0043,16'h0002,-16'h00ad,-16'h01dc,16'h00c8,16'h0071,16'h00a7,-16'h0022,-16'h0055,16'h00cb,16'h00df,-16'h008e,16'h010a,-16'h0025,16'h002a,-16'h00b4,-16'h0270,-16'h002c,16'h0047,16'h0074,-16'h0099,16'h00c1,-16'h00ae,-16'h0153,16'h013d,-16'h0037,16'h00cd,16'h0038,16'h0116,-16'h014d,-16'h002c,-16'h00b6,16'h00b9,16'h0119,-16'h0156,-16'h00bf,16'h0005,16'h0065,-16'h0122,-16'h0084,16'h000a,16'h0073,-16'h005f,16'h00dc,16'h000f,16'h005c,16'h00b4,-16'h0070,16'h0061,-16'h00f3,-16'h0072,-16'h026a,16'h0152,16'h0044,16'h007b,16'h00c1,16'h0148,16'h00f6,16'h00ab,16'h00ab,-16'h0071,16'h00a8,16'h009d,-16'h0089,16'h0001,16'h0071,-16'h0041,-16'h031f,16'h009f,16'h003d,16'h00b7,-16'h0044,-16'h005b,16'h0160,16'h0190,-16'h00e6,16'h012f,16'h002a,16'h0057,-16'h006d,-16'h02dc,16'h0091,16'h0011,16'h0053,-16'h0077,16'h0031,-16'h0080,-16'h0191,16'h008b,-16'h0035,-16'h011c,-16'h000a,16'h00da,-16'h0211,-16'h0027,-16'h0126,16'h0038,16'h0103,-16'h019d,-16'h0150,-16'h004e,-16'h0042,-16'h0129,-16'h0020,-16'h0049,16'h0001,-16'h00de,16'h00b7,16'h0026,16'h0085,16'h010a,-16'h0011,16'h007c,-16'h0060,-16'h011f,-16'h01ac,16'h0155,16'h0006,16'h0107,-16'h003c,16'h00b7,16'h01c5,16'h0171,16'h004a,16'h002c,16'h004a,16'h00fa,-16'h0083,16'h0011,-16'h0036,16'h007a,-16'h02d2,16'h0059,16'h0021,16'h00d0,-16'h0060,16'h000c,16'h0130,16'h016e,16'h002b,16'h00ef,16'h0113,-16'h0007,-16'h002c,-16'h03a5,16'h0070,-16'h003f,16'h0091,16'h0043,16'h0053,-16'h0006,-16'h0141,-16'h0096,-16'h0024,-16'h0270,16'h00b6,16'h00a0,-16'h0110,-16'h0073,-16'h004a,16'h0012,16'h00a1,-16'h017d,-16'h0079,16'h0054,-16'h01cd,-16'h007f,-16'h0077,-16'h002d,16'h007f,-16'h01ac,16'h006c,-16'h001a,16'h0004,16'h0065,16'h00aa,16'h0138,-16'h00a5,-16'h00c2,-16'h0169,16'h0161,-16'h008e,16'h015d,-16'h013f,16'h0001,16'h01bb,16'h006c,-16'h002d,-16'h009f,16'h007f,16'h010d,-16'h007b,16'h00d1,16'h008a,16'h00bb,-16'h02a7,-16'h005d,-16'h0021,16'h0035,16'h0062,16'h004e,16'h00e8,16'h014f,16'h00d3,16'h0097,16'h0009,16'h003e,-16'h000c,-16'h0351,-16'h003a,16'h0044,16'h0004,-16'h0049,16'h004f,-16'h00df,-16'h015a,-16'h0173,-16'h003c,-16'h0107,16'h010d,-16'h0003,-16'h00c1,-16'h0096,16'h00b8,-16'h004f,-16'h0016,-16'h013d,16'h008d,16'h008a,-16'h01c5,16'h0006,-16'h008a,-16'h007e,16'h006c,-16'h0179,16'h0091,-16'h01b9,16'h000a,-16'h0037,16'h01d1,16'h015a,-16'h0133,-16'h0046,-16'h015c,16'h0165,-16'h0095,16'h01fa,-16'h0188,16'h0066,16'h01d4,-16'h0042,16'h00c9,-16'h00f2,16'h00b4,16'h005f,-16'h00dc,16'h00c0,16'h00bb,16'h00d2,-16'h01f4,-16'h00e8,16'h0018,16'h0046,16'h006b,16'h006f,16'h0116,16'h018f,16'h0124,16'h006d,16'h0027,-16'h0019,-16'h0022,-16'h030c,16'h0007,16'h0056,16'h006c,16'h0000,16'h0029,-16'h014b,-16'h0233,-16'h01b5,-16'h0035,16'h0101,16'h0145,16'h0085,16'h0038,-16'h0077,16'h0075,-16'h0034,-16'h0141,-16'h00f1,16'h00f5,-16'h00dc,-16'h0195,-16'h006c,-16'h003d,-16'h00c7,16'h00a9,-16'h00f8,16'h00ca,-16'h0250,-16'h0073,-16'h0070,16'h01f2,16'h0092,-16'h0107,16'h006d,-16'h0146,16'h0137,-16'h009f,16'h01c1,-16'h0288,16'h0045,16'h01bc,-16'h0097,16'h017f,-16'h0178,16'h00e1,16'h003c,-16'h004b,16'h011c,-16'h005e,16'h0100,-16'h0236,-16'h0272,16'h0001,16'h00b1,16'h00dd,16'h0009,16'h008e,16'h01b9,16'h011c,16'h00f6,-16'h000f,-16'h00ba,-16'h002f,-16'h0312,16'h0026,16'h007e,16'h0074,16'h005f,-16'h0050,-16'h0131,-16'h01f6,-16'h0218,-16'h00d4,16'h0236,16'h00dd,16'h003f,16'h00c5,-16'h0015,16'h006b,16'h000b,-16'h01c9,16'h002c,16'h0167,-16'h017b,16'h0020,-16'h00ab,-16'h0041,-16'h00a5,16'h0034,-16'h0046,16'h00fc,-16'h0273,-16'h0062,16'h0019,16'h0076,-16'h003c,-16'h0002,16'h00c1,-16'h0128,16'h00a5,-16'h00c5,16'h00a7,-16'h0270,16'h0073,16'h011e,-16'h0046,16'h0137,-16'h01f4,16'h0019,16'h0042,16'h001a,16'h0163,-16'h00ad,16'h0113,-16'h0208,-16'h0228,16'h0018,16'h005e,16'h0074,16'h012a,16'h002f,16'h015c,16'h00bb,16'h004a,-16'h0042,-16'h0092,-16'h009a,-16'h0268,16'h006a,16'h005e,16'h008a,16'h0073,16'h0033,-16'h017f,-16'h01e3,-16'h02c7,-16'h0117,16'h01de,16'h0175,16'h003e,16'h005e,16'h005f,16'h012a,16'h0058,-16'h0129,16'h012d,16'h0064,-16'h0156,16'h0193,-16'h0114,-16'h003e,-16'h00ed,16'h0042,16'h0075,16'h00c4,-16'h00e2,-16'h005e,16'h0068,-16'h01af,-16'h0049,-16'h002b,16'h009f,-16'h00cd,16'h0096,16'h0044,-16'h0106,-16'h02cc,16'h008d,16'h0111,16'h0086,16'h0085,-16'h0254,16'h0018,16'h0045,16'h009d,16'h01c5,-16'h0029,16'h0144,-16'h0128,16'h008d,-16'h0003,16'h0052,16'h00f6,16'h008e,-16'h00b1,16'h01e2,16'h0076,16'h0001,-16'h0030,-16'h00a5,-16'h00c7,-16'h024d,16'h00ff,16'h00c3,16'h00e9,16'h007a,16'h007d,-16'h00d2,-16'h01b2,-16'h03e8,-16'h0079,16'h0049,16'h0012,16'h0095,16'h0089,-16'h0017,16'h0110,16'h00a8,-16'h008e,16'h012d,16'h0057,-16'h0194,16'h0204,-16'h00f0,-16'h008f,-16'h00f9,-16'h003c,16'h0090,16'h00b0,16'h00a0,-16'h008c,16'h00bd,-16'h0202,16'h014b,16'h0062,16'h0084,-16'h00cf,16'h0133,16'h00d6,-16'h0100,-16'h0256,16'h0109,16'h018a,16'h0056,-16'h0009,-16'h0202,-16'h000b,16'h0074,16'h0021,16'h0126,16'h0020,16'h0173,-16'h00b9,16'h0158,16'h002f,-16'h0005,16'h0091,-16'h001d,-16'h0009,16'h019e,16'h0024,-16'h001c,-16'h001b,-16'h0012,-16'h0050,-16'h0212,16'h0155,16'h00ed,16'h0141,16'h009d,16'h00e5,-16'h00e5,-16'h004d,-16'h0347,-16'h000e,-16'h0191,-16'h0181,16'h0013,16'h00ac,-16'h0028,16'h00fa,16'h0097,16'h006a,16'h00ea,16'h0069,-16'h0125,16'h0205,-16'h00bd,-16'h009b,-16'h00a7,-16'h0057,16'h0053,16'h00ce,16'h01a5,-16'h0129,16'h0175,-16'h01b5,16'h01d2,16'h0075,-16'h0127,-16'h00cf,16'h019a,16'h006f,-16'h00ca,-16'h0185,16'h0110,16'h00e2,16'h00a7,-16'h0028,-16'h01a7,16'h005a,16'h0073,16'h00a6,16'h0129,16'h002e,16'h0190,-16'h00bb,16'h015a,16'h0050,16'h0000,16'h00d8,-16'h000f,16'h001a,16'h0200,16'h00fb,16'h005d,16'h0049,-16'h00b4,-16'h001c,-16'h01e8,16'h0102,16'h0081,16'h0137,16'h0010,16'h0036,-16'h0139,-16'h002f,-16'h0146,-16'h0020,-16'h01df,-16'h0189,16'h0046,16'h008d,-16'h002e,16'h014f,16'h0122,16'h002a,16'h00b8,-16'h0031,-16'h0125,16'h017c,-16'h0111,16'h0000,-16'h00b3,-16'h002b,-16'h00cc,-16'h0022,16'h01d2,-16'h00b4,16'h00bb,16'h0005,16'h0109,16'h0078,-16'h01a0,-16'h0038,16'h00f9,16'h00dc,-16'h0117,-16'h009e,16'h00f1,16'h00db,16'h0097,-16'h0049,-16'h0224,16'h0033,16'h0096,16'h00f7,16'h006d,-16'h0007,16'h01c8,-16'h0001,16'h018f,16'h00a8,-16'h0009,16'h009f,16'h0071,16'h002b,16'h024a,16'h00bf,16'h0056,16'h0034,-16'h0085,-16'h0043,-16'h020b,16'h015a,16'h0085,16'h0125,-16'h0085,-16'h003e,-16'h00c8,-16'h000d,-16'h004f,16'h0060,-16'h00bb,-16'h0170,-16'h0041,16'h006b,-16'h00e3,16'h00eb,16'h0084,16'h000c,16'h00d6,-16'h0081,-16'h0027,16'h00cb,-16'h010e,16'h00a0,-16'h0142,16'h0149,-16'h0144,-16'h0080,16'h01f2,-16'h006f,16'h00a6,16'h0185,-16'h00e7,-16'h000c,16'h0032,-16'h0077,16'h00b9,16'h006f,-16'h00cd,16'h0035,16'h016e,-16'h0049,16'h006d,-16'h0122,-16'h0269,16'h0020,16'h0096,16'h0055,16'h0083,-16'h005c,16'h0169,16'h0039,16'h012a,16'h0057,16'h0057,16'h004a,16'h009c,-16'h0058,16'h0284,16'h0138,16'h0026,16'h007d,16'h0011,-16'h002b,-16'h01ce,16'h013f,16'h018c,16'h017e,-16'h0049,-16'h0004,-16'h00d7,16'h001f,16'h00b7,16'h009e,16'h0093,-16'h000a,-16'h0046,16'h0020,-16'h0058,16'h014a,16'h0080,16'h0052,16'h00dc,-16'h00c6,-16'h0039,16'h0007,-16'h004d,16'h00c8,-16'h014e,16'h0152,-16'h0116,-16'h0044,16'h022f,-16'h0056,-16'h00b3,16'h012a,-16'h0253,16'h0012,16'h00af,-16'h009d,16'h0045,16'h008e,-16'h0189,16'h00f1,16'h007d,16'h0030,16'h00c2,-16'h008a,-16'h01e6,16'h0020,16'h0138,16'h0076,16'h0086,-16'h0046,16'h0167,16'h0096,16'h000b,16'h0052,16'h000f,16'h00e0,16'h0048,-16'h00ce,16'h0213,16'h01d2,16'h0087,16'h0058,-16'h00cc,-16'h002d,-16'h01ad,16'h008f,16'h017d,16'h00eb,-16'h00a5,16'h003e,-16'h0146,16'h00a3,16'h00ce,16'h000c,16'h01b0,16'h00ec,-16'h0073,16'h009e,-16'h00d2,16'h00d3,16'h006d,-16'h004f,16'h00b8,-16'h00be,-16'h0095,-16'h00ed,-16'h0085,16'h008d,-16'h0129,16'h0158,-16'h00c8,-16'h004e,16'h0208,-16'h0042,-16'h0201,16'h00b7,-16'h0124,16'h0040,16'h0018,-16'h0052,-16'h0029,16'h0095,-16'h011e,16'h012b,16'h0060,-16'h0001,16'h00be,-16'h0038,-16'h00fb,-16'h00af,16'h0138,16'h0048,16'h0077,16'h0003,16'h0024,16'h00da,-16'h0066,16'h00a9,-16'h001a,16'h00f9,16'h00db,-16'h00eb,16'h01e6,16'h0126,16'h0008,16'h005d,-16'h0196,-16'h0023,-16'h0188,-16'h0008,16'h0163,16'h0128,-16'h0094,-16'h0030,-16'h009c,16'h00ed,16'h00c1,16'h001d,16'h014b,16'h00ef,-16'h0086,16'h0030,-16'h00fd,16'h0121,16'h007d,16'h001f,16'h00c1,-16'h00b8,-16'h006e,-16'h00ce,16'h001a,16'h00a0,-16'h0138,16'h0074,16'h0025,16'h0032,16'h0169,-16'h0049,-16'h0233,16'h00da,16'h00b8,16'h0088,16'h0010,-16'h0044,-16'h008f,16'h0068,-16'h0087,16'h00da,-16'h001a,16'h004a,16'h011c,16'h0033,-16'h0125,-16'h01a9,16'h00b0,16'h0003,16'h001e,16'h00e0,-16'h0081,16'h0114,-16'h00cf,16'h0046,-16'h001e,16'h00d9,16'h00a8,-16'h00b1,16'h017c,16'h00cf,16'h0045,16'h00d9,-16'h010c,16'h002b,-16'h019c,-16'h014f,16'h01c5,16'h00fb,-16'h014a,16'h00b5,16'h0077,16'h0069,16'h000a,16'h0004,16'h0102,16'h0076,-16'h0055,16'h0034,-16'h0140,16'h00bc,16'h0080,-16'h003b,-16'h0002,-16'h00b8,-16'h00c0,-16'h0031,-16'h0105,16'h0082,-16'h0131,-16'h001f,16'h00c8,16'h008e,16'h0121,-16'h0020,-16'h033a,16'h0046,16'h00da,16'h0019,16'h000c,-16'h005b,-16'h0131,-16'h0023,-16'h007a,16'h0117,16'h0000,16'h0020,16'h007d,16'h00cd,-16'h00d8,-16'h0153,16'h00d9,16'h0019,-16'h0038,16'h0048,-16'h00f6,16'h00ff,-16'h008c,16'h008a,16'h0007,16'h00ee,16'h000a,-16'h00fa,16'h011e,16'h00b9,16'h001a,16'h0123,-16'h0123,16'h000a,-16'h0198,-16'h0199,16'h0133,16'h0158,-16'h00f8,16'h0180,16'h005a,-16'h0035,-16'h00dc,-16'h003e,16'h0117,16'h00f3,-16'h009c,16'h0032,-16'h0164,16'h0138,-16'h000d,16'h0035,16'h0016,-16'h0035,-16'h010f,-16'h002b,-16'h0052,16'h001e,-16'h011a,16'h0007,16'h00d7,16'h0129,-16'h000d,-16'h0048,-16'h005a,16'h002a,16'h0154,16'h000a,-16'h0071,16'h005f,-16'h0154,-16'h003d,-16'h0090,-16'h0038,-16'h001d,-16'h010f,16'h0084,16'h007c,-16'h0117,-16'h0115,16'h010c,16'h0061,16'h0032,16'h0068,-16'h0111,16'h0068,16'h003a,16'h00ed,-16'h0043,16'h00e3,16'h0047,-16'h019f,16'h0157,-16'h0077,16'h0061,16'h0047,-16'h0110,16'h0009,-16'h0162,-16'h0178,16'h00f6,16'h00e2,-16'h009c,16'h0175,16'h00f7,16'h0054,16'h0008,-16'h0065,16'h0089,16'h005d,-16'h00d1,16'h006c,-16'h0144,16'h007b,-16'h0096,-16'h00b6,-16'h0039,-16'h0013,-16'h0128,-16'h0070,16'h0036,-16'h004c,-16'h010b,16'h0071,16'h0102,16'h0111,-16'h00b7,-16'h0019,16'h0084,-16'h001a,16'h00e7,16'h0005,-16'h0091,16'h0039,-16'h0059,16'h006c,16'h0054,-16'h0089,16'h008c,-16'h00d7,16'h00ce,16'h00cf,-16'h0092,-16'h0009,16'h008c,16'h00d2,16'h0005,16'h002b,-16'h0143,16'h006f,16'h0031,16'h0100,16'h001b,16'h00cb,16'h0045,-16'h0256,16'h00d9,-16'h014c,16'h000c,16'h008c,-16'h0221,-16'h0073,-16'h0199,-16'h01c8,16'h0071,16'h00f9,-16'h015e,16'h012d,16'h017f,16'h00dc,16'h0065,-16'h00cf,-16'h0023,-16'h010a,-16'h0093,16'h0057,-16'h014f,16'h008d,-16'h00dc,-16'h0253,-16'h0013,-16'h00c5,-16'h0120,-16'h0018,16'h00b8,16'h0019,-16'h009a,16'h00e7,16'h013e,16'h00b2,-16'h0030,-16'h008d,16'h01cd,-16'h0077,-16'h0144,-16'h0003,-16'h00d3,16'h0062,-16'h001b,16'h0005,16'h00b8,-16'h00cb,16'h007d,-16'h00eb,16'h0078,16'h00fa,-16'h006b,16'h0033,16'h0087,16'h008d,16'h0005,16'h004a,-16'h0135,16'h00c8,16'h0068,16'h00a2,16'h003a,-16'h0038,-16'h0036,-16'h01cf,16'h0047,-16'h01ff,-16'h0001,16'h009e,-16'h02e4,-16'h0018,-16'h0184,-16'h0126,16'h0101,16'h00c7,-16'h012b,16'h00c5,16'h01c7,16'h00e8,16'h00c2,-16'h0126,-16'h001c,-16'h023a,-16'h0161,16'h007a,-16'h00a7,16'h001f,-16'h00fc,-16'h042b,-16'h0120,-16'h0072,-16'h011a,16'h011e,16'h00dc,-16'h02c7,-16'h00d6,16'h00d2,16'h0132,-16'h00dd,-16'h0039,-16'h0027,16'h01d2,-16'h00f1,-16'h01fe,-16'h006f,-16'h00af,16'h0036,16'h0044,16'h009e,16'h0108,-16'h0107,16'h008d,-16'h0050,16'h004b,16'h0092,-16'h00eb,16'h0046,16'h0080,16'h0073,-16'h0002,16'h0033,-16'h0064,16'h0135,16'h0035,16'h00ce,16'h0085,-16'h0155,-16'h0086,-16'h0038,16'h004f,-16'h02e8,16'h0060,16'h0058,-16'h03a2,-16'h0065,-16'h01db,-16'h009f,16'h00ec,16'h00a3,-16'h0076,16'h0077,16'h0120,16'h012d,16'h00a8,-16'h0033,16'h001b,-16'h0371,-16'h01b2,16'h0082,-16'h0010,-16'h001f,-16'h009d,-16'h04cf,-16'h0171,16'h001b,-16'h000c,16'h0139,16'h0081,-16'h0617,-16'h012c,16'h0042,16'h00df,-16'h017f,16'h0054,16'h001b,16'h0076,-16'h00d2,-16'h0304,-16'h0066,16'h0067,16'h0091,16'h008f,16'h001c,16'h0113,-16'h005b,16'h00a2,-16'h0066,16'h00de,16'h008e,-16'h00ff,16'h0094,16'h00d1,16'h0064,16'h0034,16'h0057,-16'h00f0,16'h012c,16'h007b,16'h00b9,-16'h0010,-16'h01ae,16'h0020,16'h00cd,16'h0046,-16'h0301,-16'h0055,16'h00a6,-16'h02f1,16'h0057,-16'h023b,-16'h0057,16'h00a1,16'h0143,-16'h004d,16'h00cf,16'h00eb,16'h0084,16'h0057,-16'h0098,-16'h0010,-16'h044f,-16'h01b4,16'h0027,-16'h0007,16'h000c,-16'h00b3,-16'h03af,-16'h019b,16'h0159,-16'h00a9,16'h0037,16'h004f,-16'h0502,-16'h0105,16'h004a,16'h006a,-16'h0356,16'h011c,16'h0020,-16'h0178,-16'h0031,-16'h0229,-16'h00b3,16'h01ad,16'h0129,16'h0006,16'h0076,16'h0035,16'h0062,16'h0076,-16'h0067,16'h00da,16'h00b3,-16'h017c,-16'h0015,16'h00dc,-16'h0008,16'h001d,16'h001d,-16'h0091,16'h0162,16'h00d7,16'h0036,-16'h0068,-16'h0102,-16'h002d,16'h011f,16'h00f9,-16'h0144,16'h001f,16'h003d,-16'h0287,16'h0098,-16'h0188,-16'h0033,16'h0059,16'h00da,-16'h0008,16'h000c,16'h00d9,16'h00d7,16'h004b,-16'h001d,16'h008d,-16'h03ad,-16'h0093,16'h002b,-16'h003f,16'h00cb,-16'h0001,-16'h025f,-16'h0156,16'h00c1,-16'h00f9,-16'h006b,16'h009e,-16'h02ea,-16'h00f1,-16'h0032,-16'h029d,-16'h0357,16'h0143,-16'h0013,-16'h0447,-16'h0056,16'h0057,-16'h0050,16'h01cc,16'h0037,-16'h003e,16'h00ca,16'h007e,16'h0072,-16'h005e,-16'h0041,16'h0090,16'h015a,-16'h0084,-16'h003c,16'h0105,-16'h001c,16'h0099,16'h006f,16'h000a,16'h0063,16'h0037,16'h0097,16'h001f,-16'h0135,16'h0075,16'h0139,16'h00a8,-16'h0022,16'h00c9,-16'h002f,-16'h02ec,16'h008d,-16'h00ed,16'h00d2,16'h00ab,16'h00b2,16'h0084,-16'h00bb,16'h0097,16'h0095,16'h004d,16'h000e,-16'h0053,-16'h014a,-16'h0049,16'h00f5,-16'h0082,16'h00a7,-16'h0063,-16'h0190,-16'h008c,-16'h0003,-16'h01cc,16'h005c,16'h0127,-16'h0308,-16'h00c7,-16'h00c0,-16'h05dd,-16'h024e,16'h00b0,-16'h0075,-16'h052d,-16'h0052,16'h0156,16'h004d,16'h00b5,16'h0027,16'h00b7,16'h00a3,16'h00e6,16'h013f,16'h002b,16'h0006,16'h00da,16'h0149,-16'h0046,16'h000a,16'h0193,-16'h0012,16'h0081,16'h0063,-16'h005c,16'h0036,-16'h0040,16'h002a,-16'h0008,-16'h00e2,-16'h0059,16'h0012,16'h0081,16'h00a2,16'h013f,-16'h0105,-16'h0279,16'h0122,-16'h00f8,-16'h001f,16'h004b,-16'h0033,16'h0101,-16'h0109,16'h00d3,16'h00a6,-16'h0091,16'h00ac,16'h003f,16'h019d,-16'h00fe,16'h0194,-16'h01ba,16'h00aa,-16'h014d,-16'h006c,-16'h0133,-16'h00c4,-16'h0290,16'h0079,16'h017f,-16'h01b2,-16'h00af,-16'h0064,-16'h054d,-16'h00e7,16'h00c2,-16'h015d,-16'h03cc,-16'h0047,16'h01bb,16'h0023,16'h001e,-16'h00cc,16'h0133,16'h0154,16'h007a,16'h01bd,16'h000e,16'h0047,16'h0173,16'h015f,-16'h00ac,16'h000b,16'h012b,16'h006d,-16'h0069,16'h009b,-16'h009f,16'h0017,16'h00b7,16'h0069,16'h003f,-16'h0075,-16'h0153,-16'h0120,16'h00cd,16'h00a8,16'h021e,-16'h01b1,-16'h0316,16'h00ff,-16'h00c7,-16'h00e2,16'h0059,16'h0003,16'h0050,-16'h00a5,16'h0092,-16'h00d7,16'h00aa,-16'h0058,16'h009a,16'h029d,-16'h020e,16'h0091,-16'h038b,-16'h006a,-16'h0041,-16'h0001,-16'h016b,-16'h00cc,-16'h0246,16'h00ea,16'h017a,16'h009e,-16'h021a,16'h0010,-16'h0423,-16'h0051,16'h006d,-16'h0109,-16'h01da,16'h00ae,16'h01b6,16'h015a,-16'h0110,-16'h017e,16'h003f,16'h0223,16'h00e2,16'h0110,16'h002d,-16'h0079,16'h0206,16'h014d,16'h0010,-16'h0060,-16'h00d7,16'h0016,-16'h0155,16'h0049,-16'h015f,-16'h01c2,16'h009d,16'h022e,-16'h013e,-16'h006e,-16'h0082,-16'h02ee,16'h007e,-16'h01f1,16'h00a0,-16'h0018,16'h00cc,-16'h0180,-16'h0112,-16'h0072,-16'h0059,16'h00c3,16'h0001,16'h000c,-16'h0236,16'h0095,16'h0298,-16'h000f,16'h002a,16'h008b,16'h0144,-16'h0107,16'h003b,-16'h0171,16'h0104,16'h0011,-16'h0073,16'h002c,16'h00d6,-16'h0024,-16'h026d,-16'h01ac,16'h00c5,-16'h009e,16'h00f7,-16'h001a,16'h00a4,16'h019f,16'h00c7,16'h00f9,-16'h005b,16'h00d2,-16'h0054,-16'h01dc,16'h0231,-16'h0028,16'h0039,16'h0103,16'h0174,16'h0116,-16'h00fb,16'h0045,-16'h00ef,16'h0038,16'h00d2,-16'h006f,16'h0000,-16'h0034,-16'h026b,-16'h0291,16'h0177,16'h0078,16'h00b6,16'h00e9,-16'h00d4,16'h002a,-16'h005f,-16'h0093,16'h00d8,-16'h0033,16'h00c6,-16'h0100,-16'h00b8,16'h003c,-16'h00b6,16'h00bd,-16'h007d,16'h00a1,-16'h01d8,16'h0067,16'h0252,-16'h005e,16'h0134,16'h0079,16'h00a3,-16'h0240,-16'h000a,-16'h015d,16'h00db,-16'h0014,-16'h00f3,-16'h0135,16'h0000,-16'h0009,-16'h0235,-16'h017a,16'h005e,-16'h00b5,16'h0056,16'h00e2,16'h006c,16'h01a6,16'h0056,16'h009b,16'h0018,16'h010b,-16'h006d,-16'h0194,16'h0282,-16'h007c,16'h00aa,16'h00a8,16'h006f,16'h00ae,-16'h0052,16'h006f,-16'h0196,16'h0025,16'h0093,-16'h00a4,16'h00ad,-16'h00b9,-16'h00f2,-16'h02d3,16'h0185,16'h0001,16'h0100,16'h0012,-16'h003c,16'h00b2,16'h0067,-16'h00ac,16'h00ac,16'h0050,-16'h000f,-16'h0150,-16'h0077,16'h006d,-16'h0061,16'h00cf,-16'h0079,16'h004d,-16'h012f,-16'h00eb,16'h01e5,-16'h0114,16'h0152,16'h0029,16'h00f9,-16'h026d,-16'h0001,-16'h0219,16'h00d1,16'h010d,-16'h010d,-16'h0111,16'h001d,16'h0030,-16'h02ab,-16'h00fa,16'h00e0,16'h0031,-16'h007b,16'h00df,16'h004a,16'h0190,16'h014b,-16'h0029,16'h0070,16'h0013,-16'h001a,-16'h027d,16'h01cf,-16'h0069,16'h00bb,16'h00b5,16'h0072,16'h00e3,16'h0059,-16'h0010,-16'h00ef,-16'h0056,16'h0091,-16'h0098,16'h009a,16'h0024,-16'h00cc,-16'h0378,16'h0135,-16'h000c,16'h0097,16'h0012,-16'h001e,16'h00f4,16'h00ed,-16'h006c,16'h00d7,16'h0005,16'h003e,-16'h0049,-16'h015b,16'h00b5,-16'h0095,16'h0002,-16'h0080,16'h00e6,-16'h0100,-16'h00f3,16'h00f5,-16'h00a8,-16'h0045,-16'h000f,16'h00de,-16'h02a3,-16'h000e,-16'h028e,-16'h0002,16'h0124,-16'h0096,-16'h00b2,16'h000f,-16'h0021,-16'h02f7,-16'h00b9,16'h0052,16'h0007,-16'h013b,16'h00fb,16'h006c,16'h00ef,16'h0110,16'h0041,16'h0055,16'h0008,-16'h00dd,-16'h02ba,16'h0243,16'h0039,16'h00ad,16'h009f,16'h0070,16'h013b,16'h0067,-16'h0021,-16'h0159,16'h000d,16'h0071,-16'h002b,16'h0042,16'h003c,16'h0000,-16'h0363,16'h01cc,-16'h0056,16'h0124,-16'h0080,16'h008d,16'h0090,16'h010d,-16'h0082,16'h00c6,16'h0035,16'h0035,-16'h007f,-16'h015d,16'h007b,-16'h001e,-16'h0008,-16'h0016,16'h0094,-16'h004b,-16'h00c4,-16'h0043,-16'h0081,-16'h0168,16'h007e,-16'h0026,-16'h01e3,16'h002a,-16'h03be,-16'h004d,16'h017c,-16'h0180,-16'h0166,16'h00a1,-16'h016e,-16'h0245,-16'h00b6,16'h0091,16'h0060,-16'h01bc,16'h00b9,16'h002f,16'h0100,16'h0112,16'h00a9,16'h0116,-16'h0089,-16'h0146,-16'h0262,16'h01da,-16'h0053,16'h013b,16'h001e,-16'h004f,16'h0215,16'h0152,-16'h0068,-16'h0132,16'h0087,16'h0037,-16'h00ec,16'h00d7,16'h001a,16'h0081,-16'h0311,16'h0061,-16'h0082,16'h0069,16'h0024,16'h0094,16'h00aa,16'h011b,16'h0099,16'h00b9,16'h0112,-16'h000c,-16'h001f,-16'h026c,16'h007f,-16'h00bd,-16'h0017,-16'h002b,16'h008d,-16'h012f,-16'h0084,-16'h01c3,-16'h0006,-16'h02be,16'h013c,16'h0012,-16'h019c,-16'h00a2,-16'h0352,-16'h006a,16'h00a8,-16'h0162,-16'h0045,16'h00d8,-16'h02c9,-16'h0157,16'h0003,16'h003d,16'h008a,-16'h01f2,16'h0070,-16'h00d5,16'h00fe,16'h0044,16'h014a,16'h01e7,-16'h00c4,-16'h00b3,-16'h01e3,16'h01cb,-16'h0033,16'h014f,-16'h00c3,-16'h0073,16'h0211,16'h0111,-16'h000e,-16'h010d,16'h00c9,16'h0043,-16'h007b,16'h0075,16'h00c5,16'h0119,-16'h01ca,-16'h005f,16'h0000,-16'h0009,16'h0038,16'h00ee,16'h00a2,16'h0178,16'h0072,16'h0093,16'h000e,16'h001f,16'h007b,-16'h0258,-16'h0010,-16'h001e,-16'h006f,-16'h008d,16'h00cf,-16'h011a,-16'h0087,-16'h02bf,-16'h0010,-16'h0108,16'h0156,-16'h0052,-16'h0097,-16'h00c9,-16'h0387,-16'h0048,-16'h0058,-16'h013a,16'h0083,16'h016b,-16'h02d6,-16'h01cf,-16'h000d,16'h0063,16'h0151,-16'h0111,16'h0032,-16'h0242,16'h00f8,16'h0028,16'h0260,16'h0146,-16'h00e8,-16'h0075,-16'h0133,16'h0175,-16'h0123,16'h010b,-16'h00f6,-16'h0075,16'h0181,16'h0028,16'h001b,-16'h013c,16'h0163,16'h0015,-16'h0022,16'h00b7,16'h00cd,16'h00fd,-16'h0169,-16'h013b,16'h004d,16'h0064,16'h00da,16'h00ac,16'h0077,16'h01a2,16'h00e1,-16'h000d,-16'h0046,16'h0097,16'h008a,-16'h027f,-16'h0024,-16'h0032,16'h005e,-16'h007b,16'h0076,-16'h0177,-16'h0114,-16'h02f8,-16'h0099,16'h0131,16'h0196,16'h003b,-16'h0006,-16'h00ad,-16'h0213,-16'h002b,-16'h012d,-16'h00cc,16'h0180,-16'h003b,-16'h0101,-16'h017b,16'h003c,16'h007f,16'h0131,-16'h00c0,16'h00a5,-16'h0202,16'h0107,-16'h0048,16'h027d,16'h0056,-16'h00b7,16'h00ca,-16'h00c0,16'h00ca,-16'h0133,-16'h0009,-16'h01ca,-16'h0003,16'h0131,16'h0005,16'h00a9,-16'h018b,16'h013e,-16'h0056,16'h0038,16'h00f6,16'h0033,16'h00d8,-16'h01c7,-16'h0235,-16'h0041,16'h00ae,16'h0035,16'h00c2,16'h002f,16'h0164,16'h0063,-16'h000b,16'h000a,16'h001f,16'h0087,-16'h02bf,-16'h002d,16'h00d3,16'h0004,-16'h0005,16'h0078,-16'h0152,-16'h006b,-16'h03c3,-16'h00bc,16'h025f,16'h0115,16'h0027,16'h00a3,-16'h0126,-16'h01e0,-16'h0068,-16'h01cd,16'h0079,16'h00cf,-16'h010e,16'h00cc,-16'h011c,-16'h007d,16'h0054,16'h0051,16'h004e,16'h0077,-16'h0184,16'h0135,-16'h0043,16'h0061,-16'h00ae,-16'h0086,16'h0155,-16'h0082,16'h00d3,-16'h0100,-16'h0110,-16'h0305,16'h0010,16'h0178,-16'h0023,16'h0190,-16'h01b5,16'h001b,-16'h004d,16'h007f,16'h011c,16'h0065,16'h01b9,-16'h014f,-16'h028f,16'h0008,16'h001f,16'h001f,16'h00f6,16'h0068,16'h012b,16'h0082,16'h0000,16'h0069,16'h0031,16'h00c1,-16'h0245,-16'h0015,16'h0065,16'h002d,16'h006d,16'h00b3,-16'h00c7,-16'h0058,-16'h04af,-16'h008f,16'h011b,16'h0066,16'h002d,16'h00bb,-16'h00d8,-16'h013e,-16'h0108,-16'h00e3,16'h019c,16'h0069,-16'h01bf,16'h018f,-16'h0114,-16'h004f,16'h0048,-16'h0060,16'h0091,16'h005b,16'h0062,16'h00e8,16'h0075,-16'h019c,-16'h00a4,-16'h0071,16'h0118,-16'h003c,16'h00dc,16'h0056,-16'h0209,-16'h0438,16'h0032,16'h01d3,-16'h001e,16'h00a4,-16'h0162,16'h005d,-16'h0045,16'h00e4,16'h00f3,16'h0175,16'h0196,-16'h0158,16'h0024,16'h0029,-16'h002a,16'h0053,16'h005f,16'h0037,16'h014e,16'h000e,-16'h00a1,16'h0025,-16'h0008,16'h0073,-16'h0280,16'h00aa,16'h0118,16'h00ce,16'h00a9,16'h0117,-16'h00a3,16'h0002,-16'h048a,-16'h0085,-16'h0003,-16'h009f,16'h0048,16'h00a0,-16'h00c8,-16'h0097,-16'h008d,-16'h0024,16'h017e,16'h0053,-16'h01cb,16'h0193,-16'h010a,-16'h006e,16'h001d,-16'h0077,16'h00e8,16'h00ab,16'h0201,16'h0117,16'h013d,-16'h0231,16'h0136,-16'h0009,16'h0021,-16'h0029,16'h0024,16'h00a5,-16'h0129,-16'h0498,16'h00e7,16'h0238,16'h007b,16'h001b,-16'h01db,16'h00c1,-16'h0079,16'h00de,16'h00ee,16'h018d,16'h0175,-16'h0003,16'h0102,-16'h0090,16'h004b,16'h00e0,-16'h0074,16'h004d,16'h0173,16'h001f,-16'h0059,16'h0046,-16'h00a1,16'h00eb,-16'h0295,16'h00f3,16'h00b4,16'h00d5,16'h00c7,16'h00da,-16'h0004,16'h00bd,-16'h02ca,16'h0014,-16'h015a,-16'h01eb,-16'h001d,16'h006a,-16'h00c6,-16'h00c7,16'h0041,16'h0060,16'h00d2,16'h0008,-16'h01d2,16'h0105,-16'h00b2,-16'h0021,16'h0065,-16'h0040,16'h009a,16'h0092,16'h01de,16'h00cf,16'h00f6,-16'h0111,16'h0152,16'h004a,-16'h0174,16'h000a,-16'h0038,16'h0138,-16'h0182,-16'h039f,16'h011b,16'h0191,16'h0099,-16'h0031,-16'h0165,16'h0032,-16'h009c,16'h00fa,16'h0086,16'h0138,16'h015d,16'h0037,16'h01c9,-16'h000f,16'h0062,16'h0046,-16'h003f,16'h0045,16'h0162,16'h0014,-16'h003f,16'h0008,-16'h00ad,16'h00a8,-16'h02a2,16'h0152,16'h0091,16'h00e3,16'h000c,16'h0082,-16'h005b,16'h0108,-16'h0080,16'h0048,-16'h0146,-16'h0186,-16'h0027,16'h00ef,-16'h0049,-16'h0079,16'h007e,16'h0027,16'h0045,-16'h0012,-16'h0180,16'h007d,-16'h00d2,-16'h0079,-16'h003a,16'h0028,-16'h00da,-16'h0035,16'h0262,16'h0109,16'h011c,16'h00d8,16'h008d,16'h0025,-16'h0180,-16'h000d,-16'h0047,16'h008f,-16'h0154,-16'h03fd,16'h0159,16'h0190,16'h0000,-16'h0065,-16'h00e7,16'h0015,-16'h0026,16'h0133,16'h0077,16'h007e,16'h00df,16'h0108,16'h011a,16'h0072,16'h0044,16'h002f,-16'h001d,16'h0043,16'h018d,-16'h0006,16'h0066,16'h0004,-16'h0014,16'h005f,-16'h026b,16'h0122,16'h00f4,16'h013c,-16'h006b,16'h0050,-16'h0011,16'h00fd,16'h00b9,16'h004d,-16'h00b2,-16'h018b,16'h002d,16'h002a,-16'h0038,-16'h00d1,16'h002c,16'h006d,16'h009e,-16'h00b3,-16'h0076,-16'h0131,-16'h018b,16'h00ca,-16'h004d,16'h00ef,-16'h013e,-16'h0054,16'h01d7,16'h010e,16'h0019,16'h0160,-16'h0183,16'h000a,16'h0017,16'h0025,-16'h004d,16'h00f8,-16'h0147,-16'h0261,16'h01aa,16'h0072,-16'h006f,-16'h00cf,-16'h014b,16'h012e,-16'h002b,16'h00b6,-16'h001c,16'h0074,16'h00d6,16'h01b8,16'h00be,16'h0044,16'h003b,16'h0095,-16'h0010,-16'h0096,16'h021c,16'h0085,-16'h0016,16'h0040,16'h00b3,16'h0032,-16'h0243,16'h0178,16'h012c,16'h00bd,-16'h001c,16'h0099,-16'h0063,16'h0063,16'h00d6,16'h00c5,16'h0007,-16'h002e,16'h0036,16'h000b,-16'h004e,-16'h00c6,16'h004a,16'h008f,16'h002c,-16'h0054,-16'h0052,-16'h01d2,-16'h0175,16'h00ec,-16'h003c,16'h0179,-16'h00fe,-16'h0098,16'h01ca,16'h0144,-16'h00e2,16'h0182,-16'h020c,-16'h007a,16'h003c,-16'h000e,-16'h0091,16'h00c2,-16'h00d3,-16'h0074,16'h0107,16'h008a,16'h00ed,16'h001d,-16'h0115,16'h00c0,16'h002e,16'h0060,-16'h006e,16'h00a3,16'h007e,16'h01ef,16'h0031,16'h0048,-16'h0007,16'h0040,16'h0059,-16'h009d,16'h0274,16'h00cb,16'h0040,16'h000d,-16'h0017,16'h004e,-16'h01f6,16'h01bd,16'h00e0,16'h00b4,16'h000a,16'h009a,-16'h00ed,16'h0099,16'h0124,16'h0048,16'h00ea,16'h008f,-16'h000c,16'h0066,-16'h004e,-16'h00c2,16'h00ba,-16'h002e,-16'h001d,-16'h006c,-16'h0064,-16'h0242,-16'h00e1,16'h00c9,-16'h0038,16'h00ba,-16'h0111,-16'h00b2,16'h01ad,16'h020b,-16'h01bb,16'h0154,-16'h0130,16'h0000,-16'h0011,16'h0021,-16'h003c,16'h011a,-16'h0035,16'h009f,16'h0048,16'h00fb,16'h0087,-16'h0069,-16'h0097,16'h0059,16'h0039,16'h003e,-16'h00a2,16'h009c,-16'h009b,16'h01d9,-16'h0067,-16'h005d,-16'h0020,16'h004a,16'h00bb,-16'h0096,16'h0223,16'h00ac,16'h007f,16'h003d,-16'h00e1,16'h002f,-16'h01ce,16'h00d0,16'h0105,16'h00e7,-16'h0042,16'h00f9,-16'h0048,16'h004d,16'h00c1,16'h003a,16'h00a8,16'h010b,-16'h007f,16'h0009,-16'h0082,-16'h0059,16'h00cd,-16'h0037,16'h0049,-16'h0070,-16'h0058,-16'h00b2,-16'h00bc,16'h00c0,-16'h0093,-16'h0016,-16'h0049,-16'h0096,16'h00c9,16'h01bf,-16'h0280,16'h0156,16'h0044,-16'h000c,16'h004b,-16'h0031,-16'h0033,16'h00a8,-16'h003e,16'h01b6,16'h001c,16'h0089,16'h0054,16'h0029,16'h0001,-16'h003c,-16'h0020,-16'h001c,-16'h0039,16'h0095,-16'h00ed,16'h0111,-16'h0105,16'h0009,16'h007a,16'h0072,16'h010f,-16'h00c6,16'h0200,16'h00a2,16'h00b9,16'h009b,-16'h00a8,16'h0061,-16'h013f,16'h005b,16'h00f4,16'h008a,-16'h0093,16'h00e4,-16'h001f,16'h0014,16'h0050,16'h008a,16'h00c7,16'h00fd,-16'h0096,-16'h0001,-16'h0122,-16'h0074,16'h001a,-16'h0085,16'h002c,-16'h0007,16'h001d,-16'h0050,-16'h0173,16'h00f8,-16'h0066,-16'h0040,16'h0135,16'h002b,-16'h009c,16'h01bd,-16'h02ac,16'h0074,16'h0104,16'h0020,-16'h0055,-16'h001e,-16'h0017,16'h003c,-16'h007d,16'h01cb,-16'h0024,-16'h0019,16'h0049,16'h0045,-16'h0069,-16'h0041,-16'h000b,16'h005b,-16'h007a,16'h0053,-16'h015e,16'h0017,-16'h0084,16'h0052,16'h007f,16'h006c,16'h0072,-16'h00ee,16'h01de,-16'h0012,16'h0046,16'h00ae,-16'h00de,16'h00ba,-16'h0133,-16'h0085,16'h004c,16'h0103,-16'h0100,16'h01b0,16'h007c,-16'h002a,-16'h00c8,16'h0010,16'h00c5,16'h0109,-16'h0101,16'h0028,-16'h01a5,-16'h00ca,-16'h004e,16'h0009,16'h0057,16'h005f,-16'h006e,-16'h008d,-16'h0187,16'h0073,-16'h00b1,-16'h00d1,16'h0144,16'h007c,-16'h0113,16'h0149,16'h0020,16'h0051,16'h0155,-16'h001b,-16'h0006,16'h0034,16'h004e,-16'h0049,16'h003e,16'h015e,-16'h004e,-16'h005d,-16'h004a,-16'h000a,-16'h001d,-16'h001c,16'h002f,16'h00f1,-16'h0077,-16'h0001,-16'h00e4,-16'h000d,16'h007a,16'h00e1,16'h000b,16'h009d,-16'h0003,-16'h00e2,16'h01f7,-16'h00b3,16'h005e,-16'h0036,-16'h0112,16'h0086,-16'h008c,-16'h00e0,16'h0058,16'h015b,-16'h00bb,16'h01ff,16'h0107,16'h001c,-16'h0025,-16'h0038,16'h0090,16'h008b,-16'h009d,16'h0082,-16'h01f4,-16'h00ef,-16'h008c,-16'h00a6,16'h003d,16'h0015,-16'h0155,-16'h006b,-16'h008e,-16'h003a,-16'h00b6,-16'h0031,16'h013a,16'h0122,-16'h0102,16'h00e3,16'h01d5,16'h0017,16'h00b0,16'h003a,-16'h006f,16'h0057,16'h00c0,-16'h005c,16'h007f,16'h00ee,-16'h0013,-16'h0077,16'h0031,16'h00cd,-16'h0028,-16'h0040,16'h003a,16'h00e6,-16'h007f,16'h000c,-16'h00b7,-16'h0089,16'h0090,16'h014e,16'h0015,16'h0037,16'h0016,-16'h0155,16'h020f,-16'h01af,16'h0032,16'h0046,-16'h00fc,-16'h0005,-16'h0103,-16'h0250,16'h0032,16'h009d,-16'h00a8,16'h012b,16'h011f,16'h00b1,16'h00a1,-16'h0067,-16'h0030,-16'h00ca,-16'h0066,16'h0086,-16'h0210,-16'h00c2,-16'h0081,-16'h0115,-16'h0010,-16'h0043,-16'h0152,16'h00fd,16'h0041,-16'h018c,-16'h00e5,16'h00b3,16'h0183,16'h010b,-16'h0039,16'h006b,16'h0230,-16'h002f,-16'h00a0,-16'h0050,-16'h0166,16'h000f,16'h0064,16'h0013,16'h00f5,16'h00e9,16'h0038,-16'h005e,16'h007e,16'h0078,16'h0094,-16'h00a6,16'h005d,16'h0066,-16'h0023,16'h007a,-16'h0057,16'h0045,16'h0109,16'h0143,16'h002f,-16'h006c,-16'h0036,-16'h0043,16'h01b9,-16'h01fc,16'h0069,16'h00ae,-16'h01d9,-16'h00a1,-16'h00e9,-16'h02b8,16'h0023,16'h008a,-16'h00f9,16'h00be,16'h00dd,16'h0152,16'h009c,-16'h0057,-16'h0072,-16'h0188,-16'h00c7,16'h0086,-16'h016a,-16'h0136,-16'h00a5,-16'h02e6,-16'h0045,-16'h0061,-16'h00cb,16'h0166,16'h002b,-16'h0498,-16'h0153,16'h003b,16'h015b,16'h0053,16'h002f,16'h0044,16'h01be,-16'h0168,-16'h0214,-16'h0094,-16'h0164,16'h0085,16'h00c5,16'h0076,16'h0119,16'h0088,16'h005a,16'h001e,16'h00ec,16'h00d5,-16'h0026,16'h0012,16'h0035,16'h0014,-16'h006a,16'h0050,-16'h00aa,16'h00ef,16'h0074,16'h007e,16'h0080,-16'h014d,-16'h0071,16'h005f,16'h00fc,-16'h021e,-16'h005c,16'h0089,-16'h01d1,-16'h00a8,-16'h015c,-16'h01db,16'h00b6,16'h008f,-16'h0091,16'h00b4,16'h0129,16'h0100,16'h00da,-16'h0069,-16'h0075,-16'h028c,-16'h015f,16'h002c,-16'h00ff,-16'h0128,-16'h0146,-16'h0511,-16'h0096,16'h00b4,-16'h00cb,16'h008d,16'h0008,-16'h0788,-16'h013f,16'h004f,16'h00a0,-16'h0154,16'h011e,16'h00ef,16'h0092,-16'h008e,-16'h0300,-16'h00c0,16'h0073,16'h008d,16'h0051,16'h0075,16'h00ed,16'h00aa,16'h00ac,16'h0001,16'h0108,16'h0135,16'h006d,-16'h0020,16'h012d,16'h0032,-16'h0024,16'h0080,-16'h004c,16'h0102,16'h00cd,16'h0007,16'h000a,-16'h0115,-16'h00c8,16'h00d3,16'h01e8,-16'h0311,-16'h0088,16'h0061,-16'h0249,-16'h0050,-16'h0124,-16'h014b,-16'h002e,16'h0104,16'h0000,16'h009f,16'h003b,16'h0102,16'h00b7,-16'h0008,16'h0002,-16'h0372,-16'h0059,-16'h0102,-16'h01a6,-16'h0098,-16'h00eb,-16'h0462,-16'h00f7,16'h018a,-16'h0090,16'h0031,-16'h0052,-16'h04d6,-16'h0109,16'h005e,16'h0003,-16'h0283,16'h018b,16'h00af,-16'h01da,-16'h0035,-16'h01dc,-16'h00e8,16'h01d1,16'h0129,16'h0055,-16'h0027,16'h00d4,16'h005d,16'h0066,16'h0069,16'h0086,16'h0114,-16'h004d,-16'h0036,16'h00d5,16'h006f,16'h0017,-16'h0029,-16'h000f,16'h0130,16'h012a,16'h0029,16'h0063,-16'h00b6,-16'h00aa,16'h0153,16'h0180,-16'h024e,-16'h0062,16'h0055,-16'h0228,-16'h0011,-16'h00f8,-16'h00c9,-16'h0016,16'h0038,16'h0086,16'h00a6,16'h00e0,16'h014e,16'h0086,-16'h009b,-16'h0020,-16'h033b,-16'h0064,-16'h00b0,-16'h0148,-16'h003b,16'h0015,-16'h0324,-16'h00b4,16'h015d,-16'h00e3,-16'h0032,-16'h001a,-16'h02fd,-16'h00c9,-16'h0016,-16'h02db,-16'h02e9,16'h020a,16'h00bf,-16'h0565,-16'h0056,16'h0125,-16'h00bf,16'h0220,16'h0036,16'h0069,-16'h0032,16'h013d,16'h0037,-16'h0091,16'h0090,16'h00c1,16'h01c2,-16'h0045,-16'h00cc,16'h011a,-16'h001e,16'h004b,16'h003a,16'h0072,16'h0160,16'h00bd,16'h007f,16'h0081,-16'h018a,-16'h0137,16'h013a,16'h0196,-16'h00ce,-16'h0021,16'h000d,-16'h0240,16'h00de,-16'h0124,-16'h0039,-16'h004f,16'h0044,16'h00fe,-16'h0116,16'h0093,16'h016e,16'h0085,16'h003f,-16'h0005,-16'h013b,16'h004c,16'h009f,-16'h01a1,-16'h003f,-16'h001f,-16'h023d,-16'h0040,16'h00be,-16'h0207,16'h0033,16'h005f,-16'h024a,-16'h005f,-16'h0075,-16'h0621,-16'h01d7,16'h01be,16'h00bf,-16'h05fa,-16'h0037,16'h01b9,-16'h0035,16'h00ee,-16'h007a,16'h010b,16'h0087,16'h00b9,16'h011c,16'h00af,16'h0110,16'h0134,16'h013d,16'h0009,-16'h00a6,16'h019e,-16'h0001,16'h00ac,16'h0005,16'h0000,16'h003d,16'h00f7,16'h005a,16'h00a7,-16'h005d,-16'h0180,16'h001b,16'h019f,16'h0012,16'h0084,-16'h004d,-16'h0192,16'h00cc,-16'h00f5,-16'h0072,-16'h007c,-16'h0093,16'h00a0,-16'h01bb,16'h009c,16'h011e,16'h0077,16'h00a0,16'h0042,16'h00c5,-16'h0091,16'h013a,-16'h01e2,16'h0009,-16'h00ed,-16'h011f,-16'h00a3,-16'h007e,-16'h0278,16'h0006,16'h0130,-16'h0172,-16'h006d,-16'h0132,-16'h053a,-16'h00af,16'h0106,16'h011c,-16'h042e,-16'h0010,16'h0195,-16'h0035,-16'h000e,-16'h00bb,16'h016d,16'h0058,16'h008f,16'h0190,16'h00d0,16'h00a9,16'h00cb,16'h013f,16'h0011,-16'h0030,16'h0148,16'h005c,16'h001c,16'h0032,-16'h00c7,-16'h005c,16'h0144,16'h005b,-16'h0004,-16'h00c2,-16'h0138,-16'h0151,16'h01e2,16'h0091,16'h020c,-16'h00d9,-16'h02a2,16'h00a1,-16'h0099,-16'h0099,-16'h009e,-16'h00a3,-16'h002b,-16'h0188,16'h0037,-16'h007b,16'h0125,16'h002d,16'h00f9,16'h01e8,-16'h01b1,16'h00d4,-16'h03b0,-16'h000d,-16'h00ed,-16'h0091,-16'h01bf,-16'h00ee,-16'h0288,16'h0094,16'h0167,16'h00b9,-16'h01a1,-16'h0014,-16'h04a7,-16'h0048,16'h0055,16'h0150,-16'h01b0,16'h0081,16'h0129,16'h004e,-16'h00e4,-16'h0193,16'h00ac,16'h01ae,16'h00a2,16'h00c6,16'h00f8,-16'h0022,16'h0140,16'h011b,16'h000f,-16'h00c9,-16'h00df,16'h006d,-16'h0191,-16'h0007,-16'h019f,-16'h0153,16'h007d,16'h0261,-16'h015c,-16'h0012,-16'h0090,-16'h0329,16'h010f,-16'h01a3,16'h0081,16'h001a,16'h008c,-16'h016e,-16'h001b,-16'h00d0,-16'h00a5,16'h00ea,-16'h001f,16'h005a,-16'h029e,16'h0098,16'h02da,16'h0079,16'h00c3,16'h0086,16'h00fb,-16'h0138,-16'h0031,-16'h01a1,16'h013a,-16'h0064,-16'h001c,16'h00b3,16'h00e8,16'h0081,-16'h0307,-16'h01bc,16'h00d0,-16'h00da,16'h00ec,16'h0055,16'h0150,16'h021b,16'h0077,16'h00b4,-16'h0033,16'h00cf,16'h0043,-16'h01f4,16'h01cb,-16'h000b,16'h00ab,16'h003b,16'h011e,16'h018c,-16'h00ec,16'h0055,-16'h008c,16'h006a,16'h0007,16'h0045,16'h0059,-16'h0096,-16'h0253,-16'h029e,16'h018e,-16'h0082,16'h0046,16'h00cf,-16'h0132,-16'h011e,-16'h0002,-16'h0086,16'h0052,16'h0041,16'h00d3,-16'h00e3,16'h0007,-16'h00a3,-16'h0072,16'h00ae,16'h0023,16'h0040,-16'h02bc,-16'h0049,16'h02c7,16'h0000,16'h007c,16'h0086,16'h00b0,-16'h0289,16'h0035,-16'h01a4,16'h008f,16'h00a9,-16'h0111,-16'h00b2,16'h00fa,16'h0032,-16'h03bf,-16'h015c,16'h0056,-16'h00a0,16'h0006,16'h011e,16'h008a,16'h01d8,16'h00da,-16'h0009,16'h0022,16'h009f,-16'h00a2,-16'h01fe,16'h0272,16'h0027,16'h015b,16'h0039,16'h00fa,16'h0121,-16'h0075,16'h0076,-16'h00af,16'h00a1,16'h008d,-16'h0095,16'h0048,-16'h0087,-16'h0126,-16'h030c,16'h0122,-16'h004e,16'h0029,16'h00b2,16'h0011,-16'h00c8,16'h002d,-16'h0053,16'h00c1,16'h0064,16'h00d3,-16'h005a,16'h0097,16'h0070,-16'h0021,16'h000a,-16'h0054,16'h0081,-16'h027a,-16'h00cb,16'h0192,-16'h0005,-16'h0007,16'h0018,16'h00ed,-16'h01e9,16'h008d,-16'h02ae,16'h0070,16'h009f,-16'h00cc,-16'h0124,16'h0074,16'h005f,-16'h0473,-16'h0142,16'h009f,16'h0031,-16'h00af,16'h00a8,16'h009f,16'h016f,16'h0127,-16'h0021,16'h0008,16'h00bd,-16'h0034,-16'h0236,16'h0268,-16'h0021,16'h0149,16'h0009,16'h000f,16'h0131,-16'h003d,16'h0016,-16'h0173,16'h0096,16'h00a7,-16'h005e,16'h007a,-16'h0082,-16'h0048,-16'h0399,16'h0171,-16'h008a,16'h00c2,-16'h0048,16'h008b,-16'h0082,16'h001c,-16'h0054,16'h0069,-16'h0032,16'h0109,16'h0040,16'h00f8,16'h0038,-16'h008c,16'h0067,-16'h0054,16'h009f,-16'h01c1,-16'h0032,-16'h001b,-16'h00c9,-16'h0048,-16'h0021,16'h00af,-16'h014a,16'h0056,-16'h031c,16'h0017,16'h014a,-16'h010f,-16'h0119,16'h0088,-16'h00a5,-16'h0497,-16'h01c0,16'h006d,16'h0009,-16'h0155,16'h0114,16'h0011,16'h010e,16'h014f,16'h0045,16'h005e,-16'h000f,-16'h00b5,-16'h0204,16'h0261,-16'h0013,16'h00f5,16'h006a,-16'h0018,16'h01d3,-16'h0003,-16'h002b,-16'h023f,16'h00a0,16'h005b,-16'h0050,16'h009a,16'h009c,16'h00c6,-16'h03b0,16'h0111,-16'h006b,16'h00cd,16'h000c,16'h00e3,-16'h0079,16'h003f,16'h0069,16'h0036,16'h0044,16'h0101,16'h00d1,16'h009c,16'h00a5,-16'h00ca,-16'h000b,16'h003d,16'h007a,-16'h012a,16'h0033,-16'h00c5,-16'h008b,-16'h01da,16'h0087,-16'h0002,-16'h00e0,16'h0053,-16'h04a2,-16'h00ad,16'h0193,-16'h00c8,-16'h0107,16'h00ef,-16'h02c9,-16'h02f6,-16'h0003,16'h007d,16'h000b,-16'h0231,16'h0043,-16'h004f,16'h00ba,16'h0106,16'h0153,16'h0127,-16'h0027,-16'h0111,-16'h0194,16'h0296,16'h0006,16'h0134,16'h0036,-16'h002d,16'h0204,16'h0078,-16'h00c9,-16'h032e,16'h0075,16'h0045,-16'h002a,16'h00b2,16'h00c4,16'h00c0,-16'h024f,16'h002f,-16'h0092,16'h004f,16'h0035,16'h013c,-16'h00a5,16'h00bc,16'h00d2,16'h0043,16'h00a7,16'h0080,16'h000f,16'h006f,16'h0073,-16'h00c1,-16'h001c,16'h0085,16'h00af,-16'h0106,16'h002e,-16'h0106,-16'h004f,-16'h02f0,16'h00e4,16'h0037,-16'h00a7,16'h001a,-16'h0525,-16'h00a1,16'h00a7,-16'h0155,-16'h0044,16'h0169,-16'h03ad,-16'h0256,16'h0091,16'h00af,16'h007d,-16'h01bb,16'h0062,-16'h0163,16'h0108,16'h0099,16'h0219,16'h018b,-16'h00a4,-16'h00fc,-16'h0120,16'h0163,-16'h003b,16'h00ef,16'h0020,-16'h000f,16'h01f4,16'h0030,16'h0015,-16'h023c,16'h00c9,-16'h0020,16'h003e,16'h00ab,16'h007d,16'h0130,-16'h0150,-16'h0094,-16'h00ac,16'h0045,16'h001c,16'h0122,16'h0047,16'h014b,16'h010c,16'h001f,16'h0044,16'h009f,16'h0028,16'h006b,16'h005b,-16'h00d6,-16'h0036,16'h0079,16'h00fc,-16'h00f4,16'h0082,-16'h025a,16'h0056,-16'h00fa,16'h01b8,-16'h001b,-16'h007b,-16'h003e,-16'h052d,-16'h0001,-16'h0068,-16'h007a,16'h007e,16'h0198,-16'h0190,-16'h0210,16'h0077,16'h0112,16'h0169,-16'h0084,16'h0005,-16'h02ba,16'h0172,-16'h0095,16'h0261,16'h0141,16'h0000,-16'h00c0,-16'h00d6,16'h00e8,-16'h00cb,-16'h000c,16'h0094,16'h0005,16'h0136,-16'h000c,16'h007d,-16'h01e1,16'h00f3,-16'h0057,16'h009d,16'h00ba,16'h0010,16'h0111,-16'h009d,-16'h00b7,-16'h003e,16'h008c,16'h004b,16'h015a,16'h0016,16'h0139,16'h0124,-16'h00d8,-16'h001d,16'h00bc,16'h0091,-16'h0031,-16'h0017,-16'h0071,-16'h0010,16'h0023,16'h00b3,-16'h008e,16'h00a3,-16'h0367,16'h0049,16'h006a,16'h00f2,16'h0027,-16'h0037,-16'h0094,-16'h0548,16'h0068,-16'h0172,16'h0006,16'h0107,16'h00d8,16'h003b,-16'h01bf,16'h00fd,16'h0144,16'h0168,16'h009c,16'h009e,-16'h0273,16'h00fd,-16'h0084,16'h01d3,-16'h0036,-16'h003a,16'h00f1,-16'h0083,16'h0077,-16'h0178,-16'h00e4,16'h00bb,16'h0018,16'h0161,-16'h0024,16'h0172,-16'h01d3,16'h010f,-16'h00c9,16'h0087,16'h0004,16'h0009,16'h020b,-16'h0096,-16'h0206,-16'h001e,16'h0068,16'h00a5,16'h0070,16'h002c,16'h0116,16'h0070,-16'h00d9,16'h0010,-16'h0016,16'h0114,16'h0014,-16'h0063,-16'h0058,-16'h000d,-16'h0035,16'h0135,-16'h0064,16'h00f3,-16'h04d9,16'h004c,16'h016c,16'h0000,16'h0008,16'h001a,-16'h0099,-16'h05eb,-16'h00b3,-16'h01cd,16'h018b,16'h00a3,-16'h007b,16'h0158,-16'h0201,16'h00a2,16'h016e,16'h00dc,16'h00f6,16'h0069,-16'h012c,16'h01b1,-16'h0004,-16'h00b5,-16'h0135,-16'h003a,16'h0251,16'h000a,-16'h0039,-16'h010f,-16'h02ae,-16'h0064,16'h007f,16'h01c6,16'h001d,16'h0158,-16'h01c6,16'h0040,16'h002a,16'h00f9,16'h0092,16'h00db,16'h0219,-16'h00f0,-16'h0226,16'h0018,16'h0083,16'h0022,16'h003c,16'h0083,16'h010a,16'h0126,-16'h0079,16'h0068,16'h0031,16'h0123,-16'h006f,-16'h000c,16'h002f,-16'h0008,16'h007c,16'h00c3,16'h003f,16'h00c8,-16'h0512,16'h000c,16'h00fc,-16'h0045,16'h001f,16'h009c,-16'h00de,-16'h04c1,-16'h00cd,-16'h006a,16'h0201,16'h0067,-16'h01a0,16'h017f,-16'h025b,16'h001c,16'h0155,-16'h0071,16'h013c,16'h004c,16'h009e,16'h01af,16'h0121,-16'h0168,16'h006a,-16'h00a4,16'h0128,-16'h0015,-16'h00b7,16'h00a6,-16'h0170,-16'h01cb,16'h00ff,16'h024d,16'h000b,16'h00fe,-16'h014b,16'h0054,-16'h0046,16'h00dc,16'h0017,16'h01cc,16'h0223,16'h005a,-16'h00c3,16'h004d,16'h003e,16'h0052,16'h0061,16'h0034,16'h0107,16'h00e6,-16'h0105,16'h0043,-16'h0010,16'h0069,-16'h00a5,16'h0034,16'h0066,-16'h003a,16'h0074,16'h0126,16'h0118,16'h0156,-16'h034b,16'h0089,-16'h0033,-16'h0108,16'h001e,16'h00fe,-16'h0179,-16'h0359,-16'h00a0,16'h0076,16'h01bb,-16'h002f,-16'h0188,16'h0162,-16'h0158,-16'h0068,16'h013a,-16'h0099,16'h0163,16'h00bf,16'h01ee,16'h0159,16'h01d5,-16'h0232,16'h011c,-16'h0063,-16'h00c5,16'h007e,-16'h0110,16'h00e9,16'h0006,-16'h0277,16'h0168,16'h0238,-16'h0002,16'h00b5,-16'h017c,16'h009e,-16'h0021,16'h00d4,16'h0049,16'h017b,16'h0149,16'h00fb,16'h00c1,-16'h003d,16'h00a5,-16'h001d,16'h0024,-16'h0066,16'h0136,16'h00a8,-16'h00a7,16'h0013,-16'h0006,16'h0050,-16'h00f7,16'h0040,16'h0047,-16'h003a,16'h00e3,16'h00e6,16'h0131,16'h0179,-16'h0062,16'h00db,-16'h01b4,-16'h0133,16'h0015,16'h006f,-16'h012f,-16'h030b,16'h0009,16'h00ae,-16'h005b,16'h002d,-16'h01bf,16'h00d6,-16'h01d0,-16'h0077,16'h0150,-16'h0033,16'h008c,16'h008a,16'h0219,16'h015f,16'h00b3,-16'h00ef,16'h00ea,16'h0027,-16'h01a4,16'h008d,-16'h00f9,16'h00a2,16'h000c,-16'h0301,16'h00c5,16'h018c,-16'h0037,16'h002c,-16'h01a1,16'h00e8,-16'h0054,16'h0064,16'h000d,16'h0188,16'h0153,16'h017c,16'h015e,-16'h0070,16'h00c6,16'h0041,-16'h0022,-16'h0092,16'h0136,16'h006b,-16'h0073,-16'h0020,16'h009a,16'h008d,-16'h0147,16'h0064,16'h0020,16'h005e,16'h0037,16'h0014,16'h005a,16'h0126,16'h017b,16'h0073,-16'h0116,-16'h0176,-16'h0015,16'h0092,-16'h0137,-16'h0257,16'h002a,16'h005b,-16'h0022,16'h000a,-16'h0188,-16'h0024,-16'h01f6,-16'h0058,16'h018e,16'h00d8,-16'h00cb,16'h0000,16'h0265,16'h01d1,16'h00fa,16'h00f3,-16'h005e,16'h002a,-16'h026d,16'h008e,-16'h0118,16'h00d1,-16'h002e,-16'h03e9,16'h0119,16'h0183,-16'h00b7,-16'h0043,-16'h0132,16'h00d0,-16'h0025,16'h0060,16'h004c,16'h00e8,16'h005c,16'h01c9,16'h0137,16'h0020,16'h009b,-16'h0005,-16'h0095,-16'h00ba,16'h00ed,16'h000b,-16'h0025,-16'h0021,16'h00b1,16'h00b3,-16'h0140,16'h00f9,16'h002b,16'h009a,-16'h0042,16'h0088,16'h012c,16'h003d,16'h01fe,16'h00cb,-16'h00e3,-16'h01b3,-16'h0059,16'h0032,-16'h015d,-16'h0219,-16'h0035,16'h0006,16'h00af,-16'h0073,-16'h0109,-16'h0228,-16'h01df,16'h0097,16'h018b,16'h00db,-16'h015d,16'h0043,16'h0152,16'h0244,16'h00b8,16'h016b,-16'h013d,16'h0023,16'h0002,16'h001b,-16'h0140,16'h0084,-16'h00c8,-16'h02ec,16'h0131,16'h0099,-16'h0069,-16'h00ab,-16'h012a,16'h0102,16'h000d,16'h001f,-16'h0058,16'h0034,-16'h0076,16'h021e,16'h0123,16'h003d,16'h00aa,16'h006c,-16'h0091,-16'h010f,16'h00b5,-16'h00de,-16'h0024,-16'h0033,16'h0125,16'h001d,-16'h013d,16'h0105,16'h0063,16'h0093,16'h003e,16'h0063,16'h0053,-16'h001a,16'h0216,16'h00f3,-16'h0043,-16'h00ca,-16'h0029,-16'h0084,-16'h01a9,-16'h01de,-16'h0041,16'h00d4,16'h006f,-16'h0063,-16'h005b,-16'h021a,-16'h01cf,16'h00a5,16'h017e,16'h0148,-16'h0138,-16'h0056,16'h0114,16'h0212,-16'h008b,16'h0111,-16'h019a,-16'h000b,16'h0047,16'h0048,-16'h0160,16'h0066,16'h0011,-16'h0253,16'h00c6,16'h0112,16'h000f,16'h0041,-16'h00d1,16'h00e9,-16'h0021,-16'h0047,-16'h0010,16'h00fc,-16'h00a1,16'h01da,16'h0033,16'h000c,-16'h0008,16'h0042,16'h0073,-16'h008f,16'h0115,-16'h0048,16'h000a,-16'h0085,16'h0183,16'h00a6,-16'h0110,16'h00c7,-16'h0082,16'h0046,16'h0091,16'h0097,16'h009e,16'h0011,16'h021a,16'h0082,16'h0011,16'h0084,-16'h0010,16'h000f,-16'h018f,-16'h01e2,16'h0059,16'h0057,16'h0023,-16'h0048,16'h0018,-16'h0204,-16'h013b,16'h0125,16'h01e2,16'h0073,-16'h01c7,-16'h0114,16'h00b5,16'h0233,-16'h01d1,16'h0165,-16'h0117,-16'h001f,16'h006f,-16'h0024,-16'h00fe,16'h00be,16'h0033,-16'h0125,16'h0015,16'h0124,-16'h0018,-16'h006b,-16'h0046,16'h00d4,-16'h007c,-16'h006d,16'h001b,16'h00fd,-16'h00fb,16'h01c2,-16'h00cb,-16'h002e,-16'h002b,16'h0016,16'h0046,-16'h0084,16'h0172,-16'h0077,16'h003b,-16'h005e,16'h0085,16'h0085,-16'h0120,16'h012c,-16'h0011,16'h006b,16'h0060,16'h0097,-16'h006f,16'h003a,16'h011e,16'h00c7,16'h0088,16'h0098,16'h0037,-16'h000e,-16'h01cf,-16'h0188,16'h0044,16'h001c,-16'h0061,-16'h00a1,-16'h0010,-16'h00cf,-16'h016c,16'h0105,16'h01cc,16'h000a,-16'h00d7,-16'h00b6,-16'h0157,16'h01c6,-16'h02a6,16'h0122,16'h001d,-16'h005e,-16'h0007,16'h0007,-16'h00eb,16'h002a,16'h0045,16'h0064,-16'h000d,16'h0103,-16'h0031,16'h0010,-16'h0028,16'h00c2,-16'h0009,16'h0008,-16'h0052,16'h0070,-16'h0140,16'h00d9,-16'h025b,16'h0017,16'h0062,16'h0005,16'h00b1,-16'h0103,16'h0138,16'h0023,16'h00a2,-16'h0030,16'h00e3,16'h0041,-16'h00dd,16'h0147,16'h0069,16'h00cb,-16'h0023,16'h0071,16'h0046,-16'h009d,16'h0041,16'h0125,16'h00ac,16'h0071,-16'h004e,16'h004d,-16'h01c7,-16'h016d,16'h0029,-16'h0072,-16'h0022,16'h0048,16'h0011,-16'h0033,-16'h0127,16'h013d,16'h018b,-16'h001c,16'h00d8,16'h0058,-16'h0202,16'h01c3,-16'h0218,16'h0055,16'h0066,-16'h0089,-16'h000d,16'h0013,16'h001d,16'h0069,16'h0000,16'h0152,-16'h0074,-16'h0005,-16'h001f,16'h0003,16'h0053,16'h0067,-16'h002a,16'h006d,16'h0005,16'h0009,-16'h010b,-16'h004f,-16'h018a,16'h0071,16'h0049,16'h0006,16'h007c,-16'h010a,16'h0162,-16'h00bb,16'h00cc,-16'h002d,16'h006c,16'h0056,-16'h0093,16'h00d0,16'h007c,16'h0167,-16'h0090,16'h01cc,16'h0027,-16'h010b,-16'h007f,16'h00a0,16'h00a8,16'h002e,16'h000c,16'h00be,-16'h019b,-16'h0204,16'h0031,-16'h0074,16'h0011,16'h0040,-16'h004d,16'h000d,-16'h0195,16'h00cd,16'h00e1,-16'h00b6,16'h015e,16'h005a,-16'h01a5,16'h0175,16'h00ea,16'h002a,16'h00f1,-16'h000e,-16'h000b,16'h0057,16'h0105,-16'h0056,16'h0096,16'h0141,-16'h0030,-16'h0074,-16'h007d,-16'h0091,16'h0016,16'h003c,-16'h00bc,16'h00e4,-16'h003a,-16'h002c,-16'h00b0,-16'h00b5,-16'h00b5,16'h008c,16'h0029,16'h0044,16'h00de,-16'h00cb,16'h01bb,-16'h0110,16'h0071,-16'h0026,16'h0053,16'h008e,-16'h0019,16'h006a,16'h00d0,16'h00f5,-16'h00f6,16'h01a0,16'h0029,-16'h0029,-16'h008a,16'h003e,16'h0090,16'h0002,-16'h0060,16'h0128,-16'h01c7,-16'h0169,-16'h00cc,-16'h00ff,-16'h0002,16'h006c,-16'h00a1,16'h00a9,-16'h00cd,-16'h003f,16'h0104,-16'h0042,16'h017c,16'h00ae,-16'h0185,16'h018b,16'h0164,16'h0092,16'h0056,-16'h004a,-16'h0064,16'h008b,16'h0110,-16'h0042,16'h0026,16'h015b,-16'h0026,-16'h003b,16'h000d,-16'h0030,16'h0027,-16'h0058,-16'h0019,16'h017c,16'h0011,-16'h0047,-16'h0085,-16'h00f9,-16'h0054,16'h018b,16'h0037,-16'h0036,16'h0056,-16'h0056,16'h0177,-16'h0130,16'h004e,-16'h002b,-16'h0054,16'h0008,-16'h004f,-16'h0101,16'h0074,16'h0054,-16'h00bc,16'h0140,16'h0035,16'h0053,-16'h005e,16'h0071,-16'h0011,-16'h00be,-16'h0058,16'h0089,-16'h0217,-16'h01bf,-16'h0105,-16'h0129,-16'h0053,16'h0019,-16'h00ec,16'h011f,-16'h0032,-16'h01b7,-16'h000a,16'h004e,16'h01c0,16'h00b7,-16'h00dd,16'h015a,16'h01de,-16'h00ae,-16'h0102,-16'h0039,-16'h0108,16'h0069,16'h00ff,16'h000d,16'h0131,16'h0196,16'h0048,16'h0070,-16'h0017,16'h0064,16'h0067,-16'h00ac,16'h0052,16'h003f,16'h0046,-16'h0033,-16'h009d,-16'h0023,-16'h003a,16'h00df,16'h0063,-16'h0126,16'h004b,16'h0022,16'h00fd,-16'h0176,16'h0034,16'h0027,-16'h001a,-16'h002f,16'h0030,-16'h01e0,16'h00d6,16'h000d,-16'h0034,16'h00cc,16'h008a,16'h011e,-16'h0007,16'h0071,-16'h008b,-16'h0115,-16'h0057,16'h0024,-16'h019f,-16'h0168,-16'h00fc,-16'h018a,16'h0023,-16'h0019,-16'h0094,16'h01b5,-16'h002b,-16'h06a4,-16'h0041,16'h0053,16'h015d,16'h009b,16'h0040,16'h0170,16'h0229,-16'h01ef,-16'h01f6,-16'h00d8,-16'h009d,16'h0044,16'h007f,16'h0093,16'h00f5,16'h010b,16'h00eb,16'h0044,16'h0005,16'h00b9,16'h0085,16'h0029,16'h00bb,16'h0085,-16'h0036,16'h0069,-16'h0006,16'h0056,-16'h0066,16'h00a2,16'h0055,-16'h0157,16'h0052,16'h0040,16'h0148,-16'h0189,-16'h004d,16'h002e,-16'h006a,-16'h0063,-16'h0032,-16'h022e,16'h0076,16'h003a,16'h0003,16'h009e,16'h0026,16'h01a5,16'h0054,-16'h000b,16'h000c,-16'h01bf,-16'h0090,-16'h0010,-16'h022f,-16'h016c,-16'h012a,-16'h0423,-16'h0009,16'h00ce,-16'h0078,16'h00cf,-16'h0089,-16'h0943,-16'h0097,16'h0083,16'h00b4,-16'h00d2,16'h0111,16'h0122,16'h0036,-16'h00a8,-16'h0123,-16'h00c2,16'h0074,16'h009a,16'h0089,-16'h00b7,16'h00c9,16'h00af,16'h00ee,16'h008d,-16'h0042,16'h012c,16'h0071,16'h006e,16'h00b9,16'h0058,-16'h0035,16'h000a,16'h004a,16'h00ba,16'h0079,16'h007e,-16'h0020,-16'h0197,-16'h00b0,16'h0123,16'h0187,-16'h01b6,-16'h0082,16'h002b,-16'h0158,-16'h0048,-16'h0049,-16'h028b,-16'h0024,16'h0052,16'h00b8,16'h001c,16'h001c,16'h018d,16'h0131,16'h0008,-16'h000c,-16'h02f5,-16'h0052,-16'h008a,-16'h0215,-16'h0148,-16'h008f,-16'h04a0,16'h003b,16'h015b,-16'h0032,16'h0037,-16'h012f,-16'h04a6,-16'h004b,16'h0085,16'h004c,-16'h02ae,16'h0137,16'h013b,-16'h027b,16'h0022,-16'h0021,-16'h0114,16'h01bc,16'h00ef,16'h003f,-16'h0063,16'h00a1,16'h00a5,16'h00f4,16'h009a,16'h0074,16'h0157,16'h003d,16'h0077,16'h0146,16'h0024,-16'h0044,-16'h0035,16'h0057,16'h0102,16'h0137,16'h0044,16'h00a1,-16'h00d6,-16'h01ea,16'h01a4,16'h01ba,-16'h0260,-16'h0017,-16'h0048,-16'h018e,-16'h005d,16'h000d,-16'h0161,-16'h00b8,16'h006c,16'h0064,-16'h009c,16'h0161,16'h0185,16'h0114,-16'h0006,-16'h0048,-16'h02e9,-16'h0021,-16'h0083,-16'h01ca,-16'h0145,-16'h0006,-16'h03e3,-16'h001c,16'h0184,-16'h0127,-16'h0074,-16'h0109,-16'h02da,-16'h00d3,-16'h00cc,-16'h036d,-16'h023e,16'h01c5,16'h00ff,-16'h05a7,16'h000e,16'h00cc,-16'h00fe,16'h019d,16'h0036,16'h0067,-16'h0006,16'h009c,16'h0072,16'h006e,16'h011a,16'h00ed,16'h017e,-16'h0088,-16'h0018,16'h00f9,-16'h0002,-16'h0074,16'h0021,16'h0034,16'h00b0,16'h00db,16'h0126,16'h010d,-16'h011e,-16'h021f,16'h0155,16'h0167,-16'h01e0,-16'h0037,-16'h0019,-16'h010f,16'h0062,-16'h0088,-16'h00af,-16'h0113,-16'h007b,16'h0101,-16'h01a7,16'h0115,16'h0118,16'h0129,16'h007c,-16'h0015,-16'h0133,16'h0006,16'h0093,-16'h01eb,-16'h00bf,16'h000f,-16'h0219,-16'h00a0,-16'h006e,-16'h021f,-16'h0033,-16'h0080,-16'h02ad,-16'h006d,-16'h012d,-16'h073f,-16'h0152,16'h011c,16'h0146,-16'h0543,16'h005c,16'h0199,-16'h0070,16'h0067,-16'h0057,16'h0147,-16'h0051,16'h0059,16'h010d,16'h0121,16'h019a,16'h005d,16'h00f9,-16'h005f,16'h000f,16'h00f0,16'h001a,16'h002f,16'h0010,16'h0066,16'h0016,16'h015d,16'h0071,16'h0096,-16'h00da,-16'h0167,-16'h004a,16'h0194,-16'h00a9,16'h00c5,-16'h0009,-16'h00e9,16'h0095,-16'h00c6,-16'h0075,-16'h0183,-16'h007f,-16'h0044,-16'h025d,16'h0069,16'h0149,16'h013e,16'h00bf,16'h0094,16'h0065,-16'h0047,16'h0068,-16'h026d,-16'h0087,-16'h011d,-16'h0145,-16'h00fe,-16'h0108,-16'h02ca,-16'h003d,16'h0005,-16'h00a0,-16'h0070,-16'h010a,-16'h0601,-16'h0100,16'h004e,16'h019d,-16'h0431,16'h0111,16'h0181,-16'h0099,-16'h0034,-16'h0032,16'h017e,-16'h0067,16'h004e,16'h0117,16'h0197,16'h0108,16'h0042,16'h00ca,-16'h0039,16'h003c,16'h0110,16'h00b7,-16'h0019,-16'h0024,-16'h006d,-16'h0093,16'h013e,16'h009c,-16'h0061,-16'h004d,-16'h00e3,-16'h0175,16'h01d9,16'h0032,16'h016b,-16'h0083,-16'h01b5,16'h006e,-16'h0056,-16'h0124,-16'h00ce,-16'h00a4,-16'h0107,-16'h024d,16'h003f,-16'h0075,16'h0154,16'h0103,16'h0156,16'h00fb,-16'h0105,-16'h0017,-16'h0406,-16'h000a,-16'h00b4,-16'h00be,-16'h01f9,-16'h0123,-16'h02da,-16'h000f,16'h0093,16'h00e8,-16'h011b,-16'h0034,-16'h0472,-16'h007a,16'h0041,16'h01cb,-16'h01b5,16'h0078,16'h011d,16'h0033,-16'h009d,-16'h00dd,16'h00eb,16'h0093,16'h006b,16'h002f,16'h01f1,-16'h0061,-16'h0005,16'h0016,-16'h0061,-16'h008e,-16'h0060,16'h0073,-16'h009e,16'h000f,-16'h0103,-16'h0142,16'h007c,16'h021e,-16'h01cf,-16'h00cb,-16'h0059,-16'h03b8,16'h01d9,-16'h0215,16'h00c5,-16'h0049,16'h00cd,-16'h0070,-16'h0026,-16'h0033,-16'h0060,16'h00ca,16'h0000,16'h005a,-16'h022e,16'h00c1,16'h0234,16'h0134,16'h00f1,16'h0057,16'h0111,-16'h0104,16'h0019,-16'h0158,16'h00ac,-16'h004a,-16'h009a,16'h0167,16'h00eb,16'h0082,-16'h0308,-16'h017a,16'h0005,-16'h012e,16'h00d9,16'h015f,16'h00bf,16'h01fc,16'h0008,-16'h0001,-16'h0083,16'h0047,-16'h0043,-16'h0114,16'h0208,16'h003c,16'h0051,16'h0131,16'h00e4,16'h017e,-16'h00b5,16'h001a,-16'h003c,16'h0133,-16'h010f,16'h005e,16'h0038,-16'h0124,-16'h015e,-16'h030c,16'h00b8,-16'h00ae,16'h0057,16'h00ce,-16'h00cb,-16'h0271,-16'h00da,-16'h00f8,16'h003e,16'h004e,16'h00ed,16'h005f,16'h00f0,-16'h006f,-16'h0044,16'h00b0,-16'h003a,16'h007d,-16'h025d,-16'h0055,16'h020a,16'h0081,16'h00b2,16'h0013,16'h00f8,-16'h0113,16'h00c8,-16'h00fe,16'h0042,16'h005b,-16'h0108,-16'h007b,16'h0090,-16'h0057,-16'h047e,-16'h01db,16'h0049,-16'h0141,16'h006a,16'h0127,16'h010e,16'h01cc,16'h0135,16'h001c,16'h003a,16'h00c2,-16'h007c,-16'h00dc,16'h02e1,16'h0064,16'h00c9,16'h00d6,16'h0146,16'h0139,-16'h0087,16'h006e,-16'h002b,16'h0135,-16'h005d,-16'h008c,16'h00b0,-16'h00d9,-16'h00ee,-16'h0327,16'h00d1,-16'h00e6,16'h0018,16'h0066,-16'h006a,-16'h033f,-16'h0073,-16'h002c,16'h0018,16'h0003,16'h0151,16'h0084,16'h0173,16'h006c,-16'h00a4,16'h0000,-16'h004f,16'h008b,-16'h02f4,-16'h006a,16'h00af,16'h00a1,-16'h0065,-16'h0027,16'h0071,-16'h005b,16'h00ec,-16'h016f,-16'h001c,16'h00de,-16'h01ad,-16'h00b9,16'h0041,-16'h011b,-16'h051e,-16'h01c8,16'h0045,-16'h014d,16'h001c,16'h0165,16'h0042,16'h012c,16'h0130,16'h0045,16'h0002,16'h00cd,-16'h001b,-16'h0130,16'h02b0,16'h00a6,16'h00b0,16'h003d,16'h00dc,16'h0170,-16'h0058,16'h004f,-16'h016d,16'h009e,16'h0056,-16'h00b8,16'h0046,-16'h003f,16'h004f,-16'h0339,16'h0133,-16'h00c1,16'h003d,16'h0052,-16'h0003,-16'h031b,-16'h0080,16'h0090,16'h008b,-16'h0067,16'h01ab,16'h011e,16'h024a,16'h0057,-16'h0092,16'h007f,16'h00b1,16'h0066,-16'h020b,16'h0011,-16'h01af,16'h0074,-16'h00e7,16'h0002,-16'h0049,16'h002b,16'h0072,-16'h01e1,-16'h00d4,16'h0192,-16'h0180,-16'h00f0,16'h0086,-16'h0225,-16'h0602,-16'h015d,16'h0016,-16'h00ae,-16'h00d4,16'h0175,16'h001b,16'h0051,16'h00cd,16'h00e1,16'h00ab,16'h006f,16'h001b,-16'h00e2,16'h025c,-16'h0025,16'h003a,16'h0030,-16'h000c,16'h01eb,-16'h004b,-16'h004f,-16'h01e1,16'h00dd,16'h00a6,-16'h0021,16'h00b6,-16'h0019,16'h00c8,-16'h0350,16'h0151,-16'h0085,16'h0096,16'h001a,16'h018c,-16'h03aa,16'h0045,16'h010b,16'h0066,16'h002b,16'h018e,16'h00a6,16'h025c,16'h003e,-16'h008c,-16'h0020,16'h00c5,16'h00b5,-16'h0113,16'h0088,-16'h023b,16'h0031,-16'h01c2,16'h006c,16'h0045,16'h005d,16'h0080,-16'h02e3,-16'h0100,16'h0164,-16'h011b,-16'h00d0,16'h0158,-16'h0309,-16'h03d3,-16'h0086,16'h0099,16'h001c,-16'h0155,16'h00b8,-16'h0089,16'h002c,16'h0099,16'h0171,16'h00d5,-16'h000c,-16'h00ad,-16'h00f1,16'h01a7,16'h0032,16'h0034,16'h0029,-16'h000d,16'h0222,-16'h0045,-16'h0036,-16'h0297,16'h00f2,16'h005d,16'h00a0,16'h009f,16'h0006,16'h0098,-16'h01aa,16'h0002,-16'h00ac,16'h0000,-16'h0004,16'h01ed,-16'h037c,16'h0094,16'h00ef,16'h0097,16'h0089,16'h0107,16'h0041,16'h0206,16'h00c8,-16'h00fc,-16'h0021,16'h00c8,16'h007a,-16'h0150,16'h012e,-16'h02b3,16'h0121,-16'h0275,16'h016a,16'h0004,16'h0046,16'h0080,-16'h0351,-16'h0011,16'h007a,-16'h0189,16'h0011,16'h01f2,-16'h02e6,-16'h02b5,16'h0033,16'h0086,16'h011b,-16'h00f8,16'h008c,-16'h02c4,16'h001f,-16'h0016,16'h021f,16'h016b,-16'h0011,-16'h006b,-16'h0088,16'h0115,-16'h00b6,16'h006a,16'h0029,16'h005e,16'h01df,-16'h0026,-16'h0081,-16'h028e,16'h000a,-16'h0032,16'h00ce,16'h008b,-16'h004d,16'h010c,-16'h00ef,-16'h006d,-16'h007b,-16'h0069,-16'h0056,16'h0218,-16'h0204,16'h010c,16'h0131,16'h001b,16'h0072,16'h00cc,16'h0008,16'h024f,16'h010e,-16'h014a,16'h0027,16'h00e6,16'h005b,-16'h0085,16'h010f,-16'h029a,16'h00ea,-16'h0156,16'h0167,-16'h0038,-16'h009f,16'h007e,-16'h0385,16'h0005,-16'h0062,-16'h0082,16'h00f6,16'h01f3,-16'h0054,-16'h0221,16'h00f6,16'h00b1,16'h0167,16'h001b,16'h0060,-16'h035d,16'h007b,-16'h0126,16'h028f,16'h009b,-16'h006e,16'h005d,16'h0009,16'h00f3,-16'h0133,-16'h0062,16'h00b3,16'h00a6,16'h00e7,-16'h003b,16'h0086,-16'h021a,16'h008f,-16'h0010,16'h009b,16'h0050,-16'h0025,16'h0138,-16'h0018,-16'h011d,-16'h0085,-16'h0023,-16'h0029,16'h0202,-16'h01b4,16'h014c,16'h00fd,-16'h007d,16'h002e,16'h0037,-16'h001b,16'h027c,16'h009c,-16'h0130,-16'h004b,16'h0058,16'h0035,-16'h0034,16'h01cb,-16'h02e0,16'h0130,16'h00b5,16'h00ab,-16'h002e,16'h002f,16'h009a,-16'h039d,-16'h003d,-16'h0113,16'h00ac,16'h008c,16'h0177,16'h0187,-16'h01e8,16'h00d4,16'h00a7,16'h0158,16'h007d,16'h0080,-16'h027c,16'h008a,-16'h00b9,16'h014e,-16'h00f1,-16'h000c,16'h01a6,-16'h000a,-16'h003d,-16'h015e,-16'h0107,16'h01a5,16'h00aa,16'h00c4,16'h0090,16'h0182,-16'h01e4,16'h0008,-16'h008f,16'h0107,16'h0045,-16'h0001,16'h01b1,16'h002b,-16'h01ea,16'h00b0,16'h007f,16'h006b,16'h011e,-16'h00d2,16'h00e1,16'h0104,-16'h005f,-16'h0009,16'h0039,16'h0037,16'h0247,16'h003e,-16'h008c,-16'h0002,16'h003c,16'h009b,16'h0046,16'h0248,-16'h0399,16'h0155,16'h011a,-16'h000f,16'h0031,16'h0007,16'h0062,-16'h0449,-16'h0011,-16'h017c,16'h0147,16'h00a0,16'h0068,16'h01b4,-16'h0218,16'h009e,16'h0141,16'h002d,16'h0120,16'h0015,-16'h0093,16'h00cf,16'h00b1,-16'h0030,-16'h0151,-16'h0057,16'h0255,-16'h0043,-16'h00ca,-16'h012c,-16'h0242,16'h014a,16'h0081,16'h01b3,16'h00ba,16'h01a8,-16'h024c,16'h0047,-16'h005e,16'h013d,16'h0018,16'h0101,16'h0217,16'h00c7,-16'h019c,16'h00e6,16'h00e9,16'h0083,16'h010d,-16'h00db,16'h00be,16'h01e1,-16'h00c8,16'h0084,-16'h0015,16'h0097,16'h0277,-16'h00a3,16'h0013,-16'h0074,16'h0041,16'h0073,16'h008c,16'h01ae,-16'h036c,16'h0105,16'h006a,-16'h00b5,-16'h0004,16'h0070,16'h0007,-16'h04c7,16'h003a,-16'h0061,16'h022e,16'h0077,-16'h010c,16'h012b,-16'h0250,16'h00b0,16'h0128,-16'h011e,16'h013d,-16'h0068,16'h0143,16'h00e7,16'h0154,-16'h0177,16'h0039,-16'h011f,16'h00e7,16'h0034,-16'h0169,16'h017a,-16'h00aa,16'h008f,16'h0130,16'h0203,16'h00e7,16'h0155,-16'h01a7,-16'h0002,-16'h0092,16'h0198,-16'h0008,16'h00dc,16'h01ad,16'h019e,-16'h0086,16'h00c0,16'h00fc,16'h0040,16'h0147,-16'h017d,16'h00df,16'h01aa,-16'h008a,16'h004b,-16'h0037,16'h0034,16'h022f,-16'h00f1,16'h006b,16'h0005,16'h00b9,16'h00ef,16'h013e,16'h0125,-16'h016d,16'h008c,-16'h0081,-16'h011d,-16'h0120,16'h005c,-16'h0053,-16'h03cb,16'h0037,16'h0071,16'h0113,-16'h0080,-16'h0109,16'h00ea,-16'h01d2,16'h0035,16'h0136,-16'h00f2,16'h0175,-16'h001b,16'h01a0,16'h00d6,16'h00f8,-16'h0183,16'h00c4,-16'h00bd,-16'h00fc,16'h005c,-16'h0209,16'h012a,16'h008a,-16'h009e,16'h010f,16'h01f1,16'h0010,16'h0043,-16'h0180,16'h0078,-16'h0170,16'h00fa,-16'h007a,16'h00a7,16'h00ae,16'h025c,16'h006e,16'h00c7,16'h01bb,-16'h0066,16'h00e5,-16'h01d3,16'h00cf,16'h013e,-16'h0035,16'h0012,16'h002e,16'h005c,16'h020b,-16'h00e5,-16'h0018,16'h0024,16'h00d4,16'h00f4,16'h013d,16'h00f0,16'h0162,16'h008d,-16'h00ad,-16'h013d,-16'h0096,16'h0063,-16'h0113,-16'h033c,16'h0095,16'h0095,16'h0016,-16'h0030,-16'h0085,-16'h005f,-16'h02a5,16'h000e,16'h013f,16'h00de,16'h0063,16'h0062,16'h0252,16'h0189,16'h008b,16'h0056,16'h00a0,-16'h00c6,-16'h025c,16'h0048,-16'h01c6,16'h00e6,16'h00c2,-16'h019a,16'h0113,16'h012c,-16'h00c0,16'h00d0,-16'h01bd,16'h0108,-16'h0093,16'h0105,-16'h0029,16'h00ce,16'h0076,16'h023a,16'h017b,16'h00a1,16'h01d7,16'h001a,16'h00ce,-16'h01f9,-16'h001f,16'h012a,-16'h00ad,-16'h0039,16'h009b,-16'h0022,16'h017f,-16'h005b,-16'h0010,16'h0038,16'h00a5,16'h010a,16'h0080,16'h012b,16'h02c9,16'h00f9,-16'h014f,-16'h00b6,-16'h006e,16'h0042,-16'h010a,-16'h02fc,16'h005a,16'h0100,-16'h0036,-16'h0032,-16'h008a,-16'h01c8,-16'h022a,-16'h0058,16'h0156,16'h00d4,-16'h00aa,16'h0094,16'h0165,16'h0185,16'h00c1,16'h0118,16'h002f,-16'h0058,-16'h0270,16'h005d,-16'h01f5,16'h0078,16'h00b9,-16'h0284,16'h0110,16'h00e2,-16'h00d9,16'h0079,-16'h00f8,16'h00e4,-16'h003b,16'h010f,-16'h0078,16'h00b0,-16'h00bc,16'h0231,16'h01a0,16'h00a6,16'h0133,16'h0056,16'h0098,-16'h016c,16'h00de,16'h00a6,-16'h003e,-16'h0016,16'h00b2,-16'h005b,16'h019a,-16'h0012,-16'h003f,16'h00f3,-16'h000d,16'h0087,16'h013e,16'h0098,16'h023c,16'h00c5,-16'h00d6,-16'h00b5,-16'h0080,-16'h0034,-16'h0157,-16'h027b,-16'h0056,16'h0019,16'h00a8,-16'h00df,-16'h003c,-16'h02e3,-16'h01f7,16'h0148,16'h0146,16'h0122,-16'h0112,16'h0073,-16'h0002,16'h0125,16'h0131,16'h0154,-16'h006f,-16'h0092,16'h0015,16'h0068,-16'h0179,16'h001e,16'h0065,-16'h0149,16'h00f9,16'h0106,16'h002b,16'h00d6,-16'h00a0,16'h007a,-16'h00a7,16'h00fe,-16'h0082,16'h002f,-16'h00f2,16'h0184,16'h011f,16'h007a,16'h014e,16'h00ec,16'h00b1,-16'h00fd,16'h00f0,16'h0002,16'h004a,-16'h0070,16'h010d,16'h0049,16'h017a,16'h0004,-16'h008a,16'h009f,-16'h0003,16'h003c,16'h00fd,16'h0034,16'h026f,16'h002c,-16'h003a,-16'h004b,-16'h0068,-16'h0115,-16'h0177,-16'h0206,16'h0025,-16'h0013,16'h00de,-16'h0057,16'h0097,-16'h02dd,-16'h0157,16'h0104,16'h0188,16'h0112,-16'h012c,-16'h0037,-16'h0087,16'h0156,-16'h0031,16'h01bf,-16'h012c,-16'h008b,16'h0080,16'h00a8,-16'h01d8,-16'h000b,-16'h003a,-16'h0140,16'h0094,16'h00de,-16'h0036,16'h0066,16'h0012,16'h0069,16'h0001,16'h009a,-16'h0088,16'h0000,-16'h016b,16'h01c8,16'h0085,16'h002a,16'h00c9,16'h0084,16'h011c,-16'h0057,16'h00df,-16'h0052,16'h0076,-16'h0056,16'h017d,16'h0066,16'h00b5,16'h004d,-16'h0077,16'h0000,16'h001c,16'h00e9,16'h0049,16'h00c1,16'h022f,16'h007a,16'h003d,16'h0027,-16'h0038,-16'h00e1,-16'h017d,-16'h01cd,16'h0093,-16'h001e,16'h004f,-16'h009b,16'h0034,-16'h0156,-16'h00e0,16'h00a0,16'h01da,-16'h0028,-16'h018f,-16'h001d,-16'h01c9,16'h0173,-16'h01a8,16'h01b9,-16'h0054,-16'h0048,-16'h0041,16'h0019,-16'h01c5,16'h006a,-16'h0018,-16'h00de,16'h0064,16'h01db,-16'h0094,16'h0090,16'h0046,16'h00cb,-16'h005f,16'h0029,-16'h001b,16'h005c,-16'h0133,16'h015e,-16'h00ec,16'h0024,16'h0032,16'h004b,16'h0153,-16'h007a,16'h00cb,-16'h004a,16'h0094,-16'h0078,16'h00fe,16'h005b,16'h007c,16'h0055,-16'h00f7,16'h0017,16'h0036,16'h005f,-16'h0051,16'h004b,16'h014f,16'h00f1,16'h0071,16'h0019,-16'h002e,-16'h0040,-16'h01e8,-16'h016d,16'h0061,-16'h0048,16'h0031,-16'h00f9,-16'h0062,-16'h0081,-16'h0063,16'h016f,16'h021b,16'h0009,-16'h00f6,-16'h0032,-16'h02d9,16'h0123,-16'h0237,16'h00ec,-16'h0001,16'h002a,16'h0049,16'h0018,-16'h0171,-16'h001e,16'h009c,-16'h0048,-16'h004f,16'h010e,-16'h0085,16'h000c,-16'h0035,16'h00c8,-16'h0001,16'h0091,16'h006b,-16'h004c,-16'h00a0,16'h002a,-16'h0228,16'h007a,16'h0079,16'h0082,16'h00c7,-16'h00aa,16'h00fc,-16'h0081,16'h00da,-16'h000c,16'h0070,16'h002f,16'h0081,16'h00ec,-16'h004a,16'h00a7,-16'h0049,16'h004c,-16'h0096,-16'h0081,16'h00d5,16'h00f6,16'h009a,16'h0061,16'h003d,-16'h0020,-16'h01d7,-16'h018b,16'h0045,-16'h006f,-16'h0125,-16'h001e,-16'h0028,16'h002f,-16'h0122,16'h0135,16'h0245,-16'h0029,16'h0144,-16'h00a4,-16'h0259,16'h009c,-16'h0207,16'h0057,-16'h0023,-16'h0076,16'h0009,16'h0071,-16'h0075,-16'h0048,16'h0044,16'h00cc,-16'h0051,16'h007a,-16'h004a,16'h0007,16'h000d,16'h00b6,16'h000b,16'h00cd,16'h0027,-16'h000c,-16'h00c7,-16'h005c,-16'h013b,16'h0079,16'h008b,16'h0056,16'h00f2,-16'h0082,16'h013d,-16'h0135,16'h014b,-16'h0050,16'h003f,16'h008a,16'h00f0,16'h00b0,16'h006e,16'h00e2,-16'h0075,16'h00a9,16'h000f,-16'h0065,16'h0019,16'h0150,16'h0054,-16'h00e3,-16'h001d,16'h00a1,-16'h0177,-16'h016f,-16'h0035,-16'h0099,-16'h00c0,16'h0066,-16'h0096,16'h0079,-16'h00d3,16'h0127,16'h0268,-16'h009d,16'h012b,-16'h0008,-16'h022e,16'h011a,-16'h004a,16'h008e,16'h00a4,16'h0046,16'h00a0,16'h002b,-16'h000a,-16'h001f,16'h0019,16'h00fc,-16'h000a,-16'h0075,-16'h009b,-16'h0005,16'h006d,16'h00d7,-16'h005c,16'h011d,16'h000d,-16'h00a7,-16'h0083,-16'h00ce,16'h0009,16'h0052,16'h002a,-16'h0003,16'h0153,-16'h0054,16'h00d2,-16'h011a,16'h0087,-16'h0080,16'h007a,16'h0018,16'h0054,16'h007f,16'h007f,16'h00b4,-16'h0031,16'h00ce,16'h005d,16'h002c,-16'h005f,16'h0157,16'h0047,-16'h003c,16'h0011,16'h0122,-16'h01b0,-16'h00fb,-16'h0040,-16'h00aa,16'h0022,16'h006e,-16'h0118,16'h0136,-16'h008b,16'h001f,16'h01bf,-16'h000e,16'h0116,16'h0005,-16'h01d8,16'h0140,16'h013a,-16'h0026,-16'h0062,-16'h0068,-16'h0029,16'h0067,16'h0042,16'h0013,16'h006c,16'h018d,16'h003d,-16'h003e,-16'h0016,16'h000c,16'h0075,16'h0078,16'h0006,16'h0108,16'h0050,-16'h00b3,16'h004d,-16'h00f9,-16'h002f,16'h0103,16'h0030,-16'h006d,16'h018a,-16'h0014,16'h00e5,-16'h017e,16'h0079,-16'h0047,16'h0028,16'h0048,16'h00f7,16'h0068,16'h00a2,16'h000d,16'h002a,16'h00fa,-16'h000f,16'h0070,-16'h0144,16'h010a,-16'h007f,-16'h002b,16'h0083,16'h0008,-16'h018c,-16'h0108,-16'h0070,-16'h00df,-16'h0011,16'h0042,-16'h0071,16'h014c,16'h002a,-16'h0225,16'h0195,16'h0093,16'h01de,16'h003a,-16'h00ab,16'h015e,16'h01f4,-16'h0063,-16'h012c,-16'h00ef,-16'h00a0,16'h0093,16'h00e9,16'h0082,16'h00f2,16'h01ff,16'h000a,-16'h0003,-16'h005e,16'h0066,16'h0072,16'h0074,-16'h0068,16'h00f2,16'h0010,16'h005b,16'h0048,-16'h00d2,-16'h003e,16'h00da,16'h0061,-16'h00ef,16'h01c8,16'h00d3,16'h0141,-16'h007a,16'h0080,-16'h011b,16'h001a,16'h0009,16'h008e,16'h000a,16'h0140,16'h0022,16'h00d0,16'h01a0,16'h000a,16'h0035,-16'h00a5,16'h00e9,-16'h00aa,16'h0003,16'h0068,-16'h007c,-16'h0135,-16'h010b,-16'h011d,-16'h00e6,-16'h0015,16'h0097,-16'h008e,16'h011c,-16'h0085,-16'h082b,16'h011f,16'h0000,16'h01b9,16'h008c,16'h0097,16'h0188,16'h016f,-16'h00fc,-16'h0135,-16'h0089,-16'h007e,16'h00a2,16'h0084,16'h00b0,16'h011c,16'h017d,16'h00e1,16'h0062,-16'h005b,16'h0154,16'h0041,16'h0070,-16'h001d,16'h005e,-16'h0042,-16'h0057,16'h005d,-16'h002b,-16'h003f,16'h00e8,16'h004e,-16'h0188,16'h01d8,16'h0085,16'h0146,-16'h003d,-16'h0042,-16'h00f2,-16'h0011,16'h0005,16'h0052,-16'h003a,16'h0068,-16'h003d,16'h013a,16'h0032,16'h0009,16'h013e,16'h0035,16'h004d,-16'h0035,-16'h014d,16'h0006,-16'h0093,-16'h01b1,-16'h0111,-16'h0123,-16'h0376,16'h0027,16'h0155,-16'h0081,16'h012f,-16'h0137,-16'h09f1,16'h00d2,16'h0054,16'h013f,-16'h006a,16'h014c,16'h00c7,-16'h0005,16'h0028,-16'h002b,-16'h0035,16'h0092,16'h0000,16'h0030,-16'h000b,16'h00e1,16'h00d7,16'h00ed,16'h0094,-16'h002b,16'h00e7,16'h0070,16'h0018,16'h0073,16'h005d,-16'h003f,-16'h0038,16'h00a8,-16'h0048,16'h008d,16'h011a,-16'h0043,-16'h0114,-16'h0079,16'h00ea,16'h0121,-16'h0034,-16'h0067,-16'h0034,-16'h00a1,-16'h003a,16'h00b2,-16'h01b1,-16'h00a1,-16'h0026,16'h00f5,-16'h00ca,16'h0095,16'h01e7,16'h00e6,16'h008e,16'h002d,-16'h026d,-16'h005d,-16'h0126,-16'h021f,-16'h011f,-16'h007f,-16'h049e,16'h0061,16'h015f,-16'h0047,-16'h0036,-16'h00e7,-16'h0545,16'h009c,16'h0036,16'h007b,-16'h0200,16'h0155,16'h013f,-16'h0200,16'h00b9,-16'h002b,-16'h0028,16'h0163,16'h0059,16'h0020,16'h0011,16'h006a,16'h0109,16'h015b,16'h009a,16'h0034,16'h0126,-16'h0033,16'h004b,16'h00a8,16'h004b,-16'h0040,-16'h003c,16'h005f,16'h00a9,16'h017a,16'h00fc,16'h005c,-16'h00b0,-16'h0325,16'h0184,16'h00e5,-16'h01cc,16'h0022,-16'h002e,-16'h00d1,-16'h0063,16'h0120,-16'h0186,-16'h0127,-16'h0089,16'h0123,-16'h02f2,16'h0146,16'h01a8,16'h014a,16'h00d0,16'h003b,-16'h0121,16'h0041,-16'h0057,-16'h01ee,-16'h010d,-16'h006d,-16'h0421,16'h0060,16'h0074,-16'h01fd,-16'h011c,-16'h00cb,-16'h0345,16'h00ba,-16'h00de,-16'h0361,-16'h01f4,16'h01dd,16'h00b4,-16'h0405,16'h011d,16'h005f,-16'h0085,16'h0186,16'h0039,16'h00a1,-16'h004e,-16'h001f,16'h0123,16'h016e,16'h00e2,16'h00dd,16'h0102,-16'h00a4,-16'h0043,16'h0154,-16'h006e,-16'h0056,16'h000c,16'h0079,16'h00af,16'h00fb,16'h010d,16'h0032,-16'h00f1,-16'h0377,16'h018f,16'h00c7,-16'h0168,16'h0041,-16'h0001,-16'h00d5,-16'h00bc,16'h0052,-16'h0132,-16'h00f3,-16'h00e6,16'h0094,-16'h0346,16'h01ba,16'h0149,16'h01c6,16'h00c2,16'h009a,-16'h00e4,16'h0047,16'h008f,-16'h01ba,-16'h0102,-16'h0047,-16'h02ba,-16'h0053,-16'h014b,-16'h0283,-16'h0139,-16'h00f2,-16'h01f7,16'h00a2,-16'h009c,-16'h070e,-16'h010a,16'h00b4,16'h00e9,-16'h041b,16'h0103,16'h0140,-16'h00ae,16'h009d,-16'h0070,16'h0142,-16'h0085,-16'h0005,16'h01b5,16'h0221,16'h015a,16'h003a,16'h0119,-16'h004a,16'h0021,16'h014b,-16'h00a8,16'h0074,-16'h006e,16'h0030,-16'h006b,16'h01a3,16'h0096,16'h008e,-16'h00a6,-16'h027a,-16'h005b,16'h0178,-16'h0171,16'h005e,16'h001c,-16'h0069,-16'h00ab,-16'h002a,-16'h01bb,-16'h00ec,-16'h004f,-16'h0030,-16'h0390,16'h00cb,16'h00ca,16'h01bc,16'h0169,16'h0054,16'h0025,16'h0021,-16'h0011,-16'h01c7,-16'h00a2,-16'h002d,-16'h01a3,-16'h0103,-16'h01c4,-16'h033f,-16'h0078,-16'h0074,-16'h00dc,16'h00a6,-16'h002f,-16'h0667,-16'h0054,-16'h00c3,16'h013c,-16'h0303,16'h00e9,16'h014a,-16'h0039,16'h002e,-16'h006a,16'h0111,-16'h00c0,-16'h0004,16'h0179,16'h0240,16'h0143,-16'h0062,16'h008a,-16'h0009,16'h0014,16'h00d6,-16'h001e,-16'h0025,-16'h0073,-16'h0004,-16'h0054,16'h0158,16'h00b7,-16'h001c,-16'h00c2,-16'h00a9,-16'h01a1,16'h0118,-16'h0020,16'h0172,16'h005a,-16'h00bf,-16'h00b0,16'h0069,-16'h0143,-16'h0096,-16'h005c,-16'h0154,-16'h02f6,-16'h0039,-16'h0043,16'h018f,16'h0150,16'h0154,16'h00a1,-16'h00ad,-16'h00b5,-16'h02c9,-16'h0061,16'h0038,-16'h00a1,-16'h0210,-16'h0184,-16'h02c9,-16'h00a2,-16'h0035,16'h0090,16'h0085,-16'h0025,-16'h04db,-16'h008f,-16'h017b,16'h01e5,-16'h01bf,16'h00bd,16'h0129,16'h002d,-16'h008e,16'h0011,16'h00de,16'h00d6,16'h0037,16'h00ad,16'h022a,-16'h0042,-16'h00a3,-16'h006a,-16'h00b9,-16'h009f,16'h0044,16'h004a,-16'h00bc,16'h0037,-16'h006a,-16'h0124,16'h0037,16'h019b,-16'h00ce,-16'h00b4,-16'h001d,-16'h0346,16'h01d7,-16'h01b4,16'h0104,-16'h0070,16'h0134,16'h00a6,-16'h0003,16'h007c,16'h00a2,16'h0142,16'h008e,16'h00ed,-16'h014c,16'h0155,16'h0176,16'h0194,16'h0131,16'h0021,16'h007f,-16'h0153,16'h0082,-16'h001f,16'h00cb,16'h002b,-16'h0057,16'h018f,16'h0080,16'h0056,-16'h02e8,-16'h0191,16'h004b,-16'h016a,16'h0132,16'h0272,16'h00bf,16'h0124,16'h004e,-16'h003c,-16'h005b,16'h005c,-16'h000f,-16'h0024,16'h029d,-16'h000b,16'h0098,16'h0109,16'h00de,16'h0122,-16'h0090,16'h0076,16'h0033,16'h0109,-16'h00d3,-16'h0024,-16'h0007,-16'h00c8,-16'h00cc,-16'h02a1,16'h00bc,-16'h0056,16'h0004,16'h0074,-16'h00a8,-16'h0234,-16'h00e5,-16'h0046,16'h00df,-16'h0069,16'h0121,16'h00e4,16'h00c0,-16'h0041,16'h004d,16'h00fb,-16'h001f,16'h00c2,-16'h0204,16'h00da,16'h006e,16'h01d0,16'h0102,16'h0012,16'h0050,-16'h00a1,16'h00ed,-16'h0046,-16'h0049,16'h0021,-16'h00f0,16'h0015,16'h00a0,-16'h0078,-16'h03f1,-16'h0100,-16'h002d,-16'h01b8,16'h0133,16'h01d0,16'h0072,16'h018d,16'h0098,-16'h00c0,-16'h0099,-16'h0006,-16'h00ab,-16'h0058,16'h02cd,16'h0114,16'h0069,16'h00aa,16'h0144,16'h0140,-16'h0082,16'h0029,16'h0006,16'h0156,-16'h00fe,-16'h00b9,16'h0060,-16'h00c2,16'h008b,-16'h0282,16'h0138,-16'h0018,16'h0045,16'h005e,-16'h002d,-16'h04b2,-16'h00bc,16'h0037,16'h00c4,-16'h0006,16'h01d9,16'h00ae,16'h0144,16'h002f,-16'h0011,16'h007f,16'h0005,16'h0071,-16'h01d8,-16'h002a,-16'h00a1,16'h0190,16'h002c,-16'h0035,16'h0002,-16'h0034,16'h0110,16'h006b,-16'h0084,16'h005f,-16'h01d5,-16'h006e,16'h0159,-16'h01e0,-16'h0498,-16'h0106,16'h002a,-16'h01c1,16'h0006,16'h0139,16'h007b,16'h00bf,16'h008c,16'h0038,-16'h0073,-16'h002c,-16'h000e,-16'h0018,16'h0280,16'h007b,16'h0069,-16'h0071,16'h00f8,16'h0180,-16'h00a9,16'h006c,-16'h00bc,16'h0135,16'h0029,-16'h0043,16'h000c,-16'h0091,16'h00ee,-16'h0255,16'h0152,-16'h0051,16'h000c,16'h0079,16'h0012,-16'h0592,-16'h0084,16'h00a1,16'h0059,16'h0028,16'h01bf,16'h008d,16'h01e2,16'h003b,-16'h0091,16'h0044,16'h0089,16'h008f,-16'h019e,-16'h000a,-16'h02d8,16'h0132,-16'h018f,16'h0004,-16'h0044,16'h00a5,16'h00c1,-16'h0034,-16'h00f2,16'h00c5,-16'h01fc,-16'h0127,16'h0140,-16'h01f1,-16'h0515,-16'h0095,16'h002c,-16'h01f6,-16'h0043,16'h01c5,-16'h002d,16'h00a5,16'h0079,16'h0136,16'h0017,16'h007d,16'h001b,16'h0068,16'h01cf,16'h008e,-16'h0020,-16'h0044,16'h00f6,16'h0214,-16'h00b5,-16'h007c,-16'h0182,16'h0128,16'h0099,16'h00b9,16'h0069,-16'h0089,16'h00a1,-16'h01c6,16'h01b7,-16'h010d,16'h0046,-16'h0004,16'h014e,-16'h056d,-16'h002e,16'h0089,16'h00a9,16'h002c,16'h01c0,16'h00a2,16'h02f4,16'h0011,-16'h014d,16'h0043,16'h00d2,16'h0080,-16'h0139,16'h00b5,-16'h03e0,16'h0140,-16'h01c3,16'h00ae,-16'h005f,16'h0096,16'h00d1,-16'h0095,-16'h0065,16'h00ee,-16'h01e9,-16'h0105,16'h0297,-16'h024c,-16'h042f,-16'h0024,16'h004d,-16'h0061,-16'h00ac,16'h00f8,-16'h00ae,-16'h0008,-16'h006b,16'h0208,16'h0097,-16'h000c,16'h0007,16'h00c9,16'h0085,16'h002a,-16'h0060,-16'h0008,16'h00f4,16'h01bc,-16'h012b,-16'h0021,-16'h0164,16'h005e,16'h0020,16'h0203,16'h0010,-16'h00b9,16'h0085,-16'h00f6,16'h00f2,-16'h00c3,-16'h007b,-16'h0055,16'h0167,-16'h063d,16'h0017,16'h006d,16'h007f,16'h0021,16'h010a,16'h0010,16'h0271,16'h0030,-16'h010d,-16'h000a,16'h01b8,16'h0023,-16'h00dd,16'h00fb,-16'h03ba,16'h018d,-16'h01c7,16'h0084,-16'h000f,-16'h0040,16'h00f0,-16'h0034,-16'h0048,16'h011f,-16'h011a,-16'h0009,16'h029d,-16'h014d,-16'h029d,-16'h000d,16'h0079,16'h006a,-16'h001a,16'h00d5,-16'h0211,-16'h0070,-16'h0107,16'h0204,16'h00cf,-16'h0010,-16'h002a,16'h00c8,16'h0082,-16'h0081,16'h0002,16'h0000,16'h00bd,16'h0120,-16'h00f6,-16'h006f,-16'h011b,16'h0070,16'h0028,16'h0239,16'h00a5,-16'h0109,16'h00ea,16'h002f,16'h001e,16'h0011,-16'h00eb,-16'h00c6,16'h01fa,-16'h069e,16'h0049,16'h009a,16'h0019,-16'h0007,16'h00d2,16'h000a,16'h029f,16'h006d,-16'h0118,16'h002c,16'h00e5,16'h009b,-16'h0148,16'h012b,-16'h0392,16'h01a5,-16'h00e5,16'h0144,16'h001c,-16'h004a,16'h0083,16'h0068,-16'h0058,16'h0085,-16'h006a,-16'h0016,16'h02ad,16'h0115,-16'h0273,16'h004b,16'h0092,16'h00fb,16'h00a2,16'h0117,-16'h026a,16'h004e,-16'h0128,16'h0236,16'h0083,-16'h000a,16'h0081,16'h0051,16'h0050,-16'h00c3,-16'h007d,16'h0071,16'h0142,16'h0172,-16'h00ff,16'h0070,-16'h00fa,16'h005d,-16'h004b,16'h0171,-16'h0027,-16'h00d3,16'h0128,16'h0063,-16'h0086,-16'h0009,-16'h00c3,-16'h0054,16'h0291,-16'h05b8,16'h004a,16'h0164,16'h000f,16'h0064,16'h00c1,16'h0022,16'h0304,16'h006b,-16'h0132,16'h0042,16'h0124,16'h008a,-16'h00d2,16'h0108,-16'h0304,16'h01df,16'h009b,16'h00ea,16'h0021,-16'h0049,16'h010e,16'h0060,-16'h00a6,-16'h00a5,16'h00ef,16'h0068,16'h0218,16'h01dd,-16'h0289,16'h00c4,16'h00e4,16'h0000,16'h0103,16'h00c1,-16'h01b8,16'h004a,16'h001c,16'h0047,-16'h00b5,-16'h002f,16'h0160,16'h0023,-16'h0049,-16'h016b,-16'h0174,16'h0104,16'h0100,16'h0137,-16'h0028,16'h0122,-16'h012c,16'h008b,-16'h0085,16'h01a3,-16'h0022,-16'h009e,16'h0206,16'h0054,-16'h0124,16'h00b8,-16'h0060,16'h0044,16'h021c,-16'h0576,16'h0099,16'h016c,-16'h005e,16'h001c,-16'h0024,16'h00ac,16'h02b6,-16'h0023,-16'h00e8,-16'h004d,16'h00e4,16'h00ac,16'h0003,16'h01f1,-16'h029f,16'h01bc,16'h0096,16'h0084,-16'h003c,-16'h00a5,16'h0110,-16'h0034,-16'h0060,-16'h00e5,16'h01a6,16'h0086,16'h011d,16'h016b,-16'h025d,16'h0135,16'h011d,-16'h01f6,16'h0105,16'h00c1,16'h0116,16'h00a7,16'h00ef,-16'h00a0,-16'h00fb,16'h002d,16'h0257,-16'h000a,-16'h00d4,-16'h0070,-16'h01cc,16'h0182,16'h0165,16'h01b7,16'h007c,16'h0142,-16'h00c7,16'h002b,-16'h0081,16'h0156,-16'h00b8,16'h0075,16'h01c5,16'h0189,-16'h0202,16'h00fc,16'h0045,16'h00d8,16'h0230,-16'h050c,16'h0080,16'h0113,-16'h000b,16'h0033,-16'h00ac,16'h006a,16'h026f,-16'h00a8,-16'h0089,16'h0032,16'h0133,16'h00c3,16'h0037,16'h0166,-16'h01cf,16'h0134,16'h0093,16'h0060,-16'h00c5,-16'h0072,16'h0137,16'h0077,16'h0015,-16'h005e,16'h019b,16'h0048,16'h0069,16'h00f8,-16'h01ff,16'h0098,16'h01a0,-16'h02da,16'h00e2,-16'h0053,16'h01dd,16'h00d0,16'h010a,-16'h0175,16'h008d,-16'h000d,16'h00e9,-16'h0039,-16'h00ca,16'h01c7,-16'h00a7,16'h0155,16'h0185,16'h0264,16'h0194,16'h0106,-16'h00fa,16'h008a,-16'h0148,16'h01be,-16'h009b,16'h000b,16'h00c4,16'h01bc,-16'h0090,16'h0195,16'h00f1,16'h00b8,16'h0276,-16'h03b9,16'h00dd,16'h0149,16'h001f,16'h0037,-16'h0071,16'h006c,16'h01c3,-16'h0138,-16'h0080,-16'h0078,16'h00ec,16'h013d,16'h00f0,16'h00bc,16'h003e,16'h012a,-16'h0043,16'h0001,-16'h0086,-16'h0090,16'h0180,-16'h000f,16'h00b1,16'h0084,16'h016f,16'h0072,16'h0008,-16'h0018,-16'h0216,16'h0075,16'h011f,-16'h0121,16'h00eb,-16'h0077,16'h01e2,16'h0114,16'h0133,-16'h00bd,16'h0119,-16'h006d,-16'h0122,16'h0042,-16'h012e,16'h0159,16'h00b7,16'h00b6,16'h01a5,16'h0172,16'h0139,16'h005a,-16'h0128,16'h00a0,-16'h013e,16'h0203,-16'h0044,16'h0003,16'h005c,16'h0203,16'h00f4,16'h0133,16'h01c6,16'h0073,16'h0279,-16'h02b9,16'h0062,16'h0165,-16'h002f,16'h0038,-16'h0041,-16'h0020,16'h021c,-16'h0105,-16'h00a0,16'h008a,16'h00b9,16'h010a,16'h00a8,16'h00dc,16'h0217,16'h011b,-16'h00b1,-16'h0056,-16'h0053,-16'h009b,16'h013a,-16'h0088,16'h0079,16'h00f0,16'h005d,-16'h001b,16'h00ce,-16'h0163,-16'h0244,16'h0082,16'h0138,16'h009d,16'h0053,-16'h0023,16'h0261,16'h00be,16'h00ac,16'h007f,16'h0001,-16'h008a,-16'h01f7,-16'h0053,-16'h0127,16'h00f8,16'h011e,-16'h004b,16'h013d,16'h00f8,16'h00bc,16'h006c,-16'h00e2,16'h012b,-16'h00b4,16'h0135,16'h0000,-16'h002d,16'h0013,16'h01d6,16'h0188,16'h0159,16'h0172,16'h00a2,16'h020a,-16'h0228,16'h008f,16'h017f,16'h0021,16'h0043,16'h0094,-16'h00a1,16'h025e,-16'h00db,-16'h00aa,16'h00e9,16'h00a2,16'h0026,16'h0100,16'h00c2,16'h025f,16'h00ea,-16'h0124,-16'h0066,-16'h0070,-16'h00d1,16'h012a,-16'h00d8,-16'h001f,16'h015d,16'h006d,-16'h000d,16'h0069,-16'h0286,-16'h0256,-16'h006d,16'h012c,16'h0094,-16'h0061,16'h0042,16'h00a8,16'h0084,16'h0130,16'h01aa,-16'h00b6,-16'h0042,-16'h019b,16'h003b,-16'h00bc,16'h00e1,16'h0196,-16'h00cc,16'h00cc,16'h0116,16'h007d,16'h00b6,-16'h00ed,16'h0062,-16'h00c2,16'h010b,-16'h002a,-16'h001c,-16'h008d,16'h01c4,16'h025b,16'h0159,16'h0171,16'h00d1,16'h01ab,-16'h00d2,16'h00b2,16'h0187,16'h0026,16'h0055,16'h0047,-16'h00a8,16'h01df,-16'h0001,-16'h00c8,16'h00da,-16'h0072,-16'h0007,16'h00c3,16'h0021,16'h020f,16'h00da,-16'h0076,-16'h0070,-16'h00ca,-16'h00c8,16'h009e,-16'h0120,-16'h0010,16'h00c2,16'h0080,-16'h007f,16'h0071,-16'h02a3,-16'h015b,16'h00d9,16'h0146,16'h003b,-16'h00c8,16'h00ca,-16'h009d,16'h0095,16'h0103,16'h01be,-16'h006f,-16'h006c,16'h00a0,16'h00b1,-16'h016a,-16'h0004,16'h0079,16'h006c,16'h0155,16'h018b,16'h00cc,16'h00bb,-16'h006e,16'h00ef,-16'h0095,16'h00e8,-16'h004a,-16'h0064,-16'h00c7,16'h01d6,16'h01b6,16'h0116,16'h0147,16'h00d4,16'h022a,-16'h0059,16'h00e7,16'h0080,16'h002b,16'h0015,16'h00a4,16'h0037,16'h0173,-16'h0079,-16'h00b2,16'h0097,-16'h00d9,16'h0019,16'h00b4,16'h009a,16'h020f,16'h00ca,-16'h002b,16'h0017,-16'h006a,-16'h0150,16'h00f3,-16'h00a4,16'h003e,16'h006b,16'h00b3,-16'h0074,16'h00bd,-16'h0267,-16'h00b3,16'h0124,16'h00b2,16'h0021,-16'h0188,16'h00b7,-16'h01df,16'h00e5,16'h0016,16'h018f,-16'h00ed,-16'h0056,16'h008a,16'h0112,-16'h0197,16'h009a,16'h0008,16'h007b,16'h0073,16'h0147,16'h0034,16'h0084,16'h004c,16'h007e,-16'h007e,16'h00c5,-16'h0038,-16'h00b1,-16'h00e4,16'h0160,16'h005c,16'h00a7,16'h0148,16'h00f1,16'h020e,-16'h000c,16'h00c9,-16'h001b,16'h0087,-16'h001f,16'h00fc,16'h0070,16'h019d,-16'h0048,-16'h00da,16'h0069,-16'h007c,16'h0027,16'h0009,16'h0123,16'h01bb,16'h0179,16'h0054,16'h00a5,-16'h00a6,-16'h0167,16'h00de,-16'h0130,16'h0039,16'h005f,16'h0050,16'h0013,16'h00c1,-16'h01d4,-16'h0017,16'h00e4,16'h011f,-16'h00ac,-16'h01e2,16'h0082,-16'h01d9,16'h00d1,-16'h00d9,16'h009d,-16'h0092,16'h0016,16'h00c9,16'h00cd,-16'h016b,16'h00d3,16'h003c,16'h00be,16'h0057,16'h0198,16'h002d,16'h0086,16'h0006,16'h0074,-16'h003e,16'h009d,16'h000e,-16'h0011,-16'h00eb,16'h014f,-16'h00d6,16'h00d4,16'h00ef,16'h00a9,16'h01ea,16'h003a,16'h00e6,-16'h0046,16'h00b3,16'h0064,16'h010f,16'h007a,16'h0139,16'h0081,-16'h013f,16'h0055,16'h0023,16'h001c,-16'h00fb,16'h011c,16'h0153,16'h0190,16'h004a,16'h0082,16'h000e,-16'h00aa,16'h00a4,-16'h00a5,16'h0080,16'h0030,-16'h005a,-16'h0086,-16'h004c,-16'h0090,-16'h004d,16'h01b3,16'h0163,-16'h0093,-16'h00f1,-16'h0048,-16'h0237,16'h010e,-16'h0199,16'h0076,-16'h0093,16'h0049,16'h00a6,16'h0098,-16'h013a,16'h0068,-16'h000b,16'h00a2,16'h0021,16'h00fb,16'h0037,16'h0098,16'h002d,16'h00cd,-16'h0062,16'h0134,16'h0061,-16'h0063,-16'h008b,16'h00af,-16'h026b,16'h013a,16'h0194,16'h006a,16'h010c,-16'h000f,16'h019e,-16'h009c,16'h0183,-16'h000e,16'h00a0,16'h003d,16'h012a,16'h0068,-16'h0041,16'h009d,16'h003a,16'h0030,-16'h0066,16'h0001,16'h0114,16'h0173,16'h0023,-16'h0017,-16'h000a,-16'h0095,16'h012f,-16'h00a3,16'h0010,16'h005c,-16'h00e4,-16'h0051,-16'h00ea,16'h0092,-16'h00a8,16'h0181,16'h01bd,-16'h010b,16'h0165,-16'h014a,-16'h0215,16'h00b4,-16'h01a6,16'h0001,16'h0022,16'h003a,-16'h0044,-16'h001c,-16'h00bf,16'h000d,16'h003f,16'h00b9,-16'h0022,16'h00fe,-16'h0004,-16'h004d,16'h0096,16'h00c3,-16'h006f,16'h01c7,16'h002d,-16'h00ab,-16'h00bf,-16'h006c,-16'h012d,16'h018c,16'h00a1,-16'h0009,16'h0167,-16'h006d,16'h0144,-16'h0117,16'h00ff,16'h000e,16'h00a2,16'h0020,16'h00f0,16'h0087,16'h0009,16'h00e9,-16'h0021,16'h0047,-16'h0001,16'h0017,16'h0010,16'h0114,16'h006e,-16'h0035,-16'h000e,-16'h0020,16'h0041,-16'h008a,-16'h0048,-16'h0048,-16'h00f4,16'h0062,-16'h00cd,16'h0137,-16'h0079,16'h0180,16'h01e6,-16'h0090,16'h013d,-16'h00cc,-16'h0186,16'h00b9,16'h0037,-16'h0053,16'h0096,16'h0084,-16'h0069,16'h0007,-16'h0028,16'h0002,16'h0110,16'h00df,16'h00c3,-16'h0015,-16'h0012,-16'h005f,16'h00bf,16'h0091,-16'h0025,16'h014e,16'h0021,-16'h014f,-16'h0030,-16'h004f,16'h00f4,16'h014d,16'h00a6,-16'h004d,16'h01f3,-16'h0042,16'h00ec,-16'h015f,16'h00d8,-16'h0019,16'h0063,16'h0073,16'h0146,16'h004c,16'h00ec,16'h00a9,16'h0086,16'h00bb,16'h003a,16'h0025,-16'h0050,16'h0170,-16'h0063,-16'h00a5,16'h0021,-16'h0026,-16'h0014,-16'h0063,-16'h0097,16'h0000,16'h000a,16'h0060,-16'h0140,16'h0141,-16'h00df,16'h0079,16'h01b2,16'h0041,16'h0186,-16'h00da,-16'h0132,16'h00fd,16'h013d,-16'h0029,-16'h0083,-16'h0042,-16'h0065,16'h0011,16'h005c,16'h000d,16'h00cd,16'h0174,16'h0017,16'h0052,16'h000c,-16'h0028,16'h006a,16'h0073,-16'h0033,16'h010c,16'h0017,-16'h0108,16'h000a,-16'h007d,16'h00d5,16'h0165,16'h0087,-16'h009d,16'h01c7,-16'h0084,16'h00fe,-16'h0157,16'h0077,-16'h0038,-16'h0071,16'h00a9,16'h0117,16'h00b7,16'h012b,-16'h0052,16'h008c,16'h0098,-16'h00b4,16'h008e,-16'h0145,16'h00fe,-16'h0028,-16'h000e,16'h006d,-16'h00ca,-16'h0055,-16'h007c,-16'h00cc,16'h00a2,-16'h002c,16'h00a2,-16'h00d5,16'h0137,-16'h005c,-16'h02d8,16'h0185,-16'h00a2,16'h01ea,-16'h00a8,16'h0022,16'h013e,16'h01e7,-16'h0013,-16'h0126,-16'h0096,-16'h00ba,16'h0055,16'h0095,16'h0068,16'h011e,16'h0181,16'h0020,16'h0033,-16'h0045,-16'h001c,16'h003e,16'h009d,-16'h004d,16'h00bb,-16'h007f,-16'h007c,16'h0089,-16'h00da,16'h000a,16'h0136,16'h0062,-16'h0094,16'h023d,16'h0048,16'h00e1,-16'h00f6,16'h00c4,-16'h0106,-16'h00af,16'h00e5,16'h00e8,16'h006f,16'h015f,-16'h0074,16'h0108,16'h0049,-16'h0019,16'h00f9,-16'h00e4,16'h0121,-16'h0039,16'h00a0,16'h006d,-16'h0121,-16'h0073,-16'h00c9,-16'h00c0,16'h0014,16'h0006,16'h01b1,-16'h0048,16'h00f2,-16'h00b3,-16'h0870,16'h015e,-16'h0051,16'h00f8,-16'h0049,16'h0125,16'h00cd,16'h0075,-16'h005d,-16'h00b4,-16'h0092,-16'h001c,16'h008e,16'h005b,16'h0105,16'h015e,16'h019f,16'h007c,16'h003a,-16'h00fa,16'h006b,16'h002e,16'h0078,16'h0012,16'h0110,-16'h0055,-16'h0050,16'h0027,-16'h0045,16'h004b,16'h0156,16'h002e,-16'h0077,16'h01e3,16'h0133,16'h00b9,-16'h0003,16'h00dc,-16'h0072,-16'h00b4,16'h0030,16'h0053,-16'h0015,16'h0066,-16'h00a6,16'h008d,-16'h00b0,16'h004c,16'h015c,16'h001a,16'h00e1,-16'h0050,-16'h00c1,16'h0035,-16'h008b,-16'h00c3,-16'h0091,-16'h00d3,-16'h020c,16'h00b4,16'h018b,-16'h00c4,16'h008e,-16'h016c,-16'h0a13,16'h0157,-16'h0068,16'h011b,-16'h00b1,16'h017a,16'h009a,-16'h0036,16'h00e0,-16'h0051,-16'h0069,16'h008d,16'h0044,16'h0042,16'h0092,16'h012f,16'h0196,16'h018c,16'h0059,-16'h00c8,16'h00a7,16'h0085,16'h0020,16'h0000,16'h00db,-16'h00c1,-16'h009c,16'h0034,-16'h0079,16'h00ef,16'h014f,16'h0000,-16'h0043,-16'h00b6,16'h006c,16'h0111,16'h0005,16'h00d9,-16'h009a,-16'h00be,-16'h0066,16'h00c3,-16'h008b,-16'h00f7,-16'h008c,16'h012f,-16'h037a,16'h00db,16'h0145,16'h0147,16'h0149,16'h0037,-16'h00cf,16'h0014,-16'h00c5,-16'h006b,-16'h00ad,-16'h0079,-16'h036f,16'h012a,16'h0100,-16'h0161,-16'h0052,-16'h01fd,-16'h055e,16'h011a,-16'h003e,16'h001b,-16'h0144,16'h017f,16'h0095,-16'h020c,16'h0130,-16'h0032,-16'h0036,16'h013d,16'h000a,16'h0045,-16'h0019,16'h000a,16'h0150,16'h0170,16'h0056,-16'h0036,16'h00be,-16'h0047,16'h0031,16'h002b,16'h005a,-16'h0058,-16'h0074,16'h00ff,-16'h0076,16'h0171,16'h01a5,16'h0014,-16'h006f,-16'h04e9,16'h00f7,16'h00ab,-16'h012d,-16'h000d,-16'h0044,-16'h00f4,-16'h00dc,16'h00dd,-16'h00e8,-16'h016a,-16'h00d2,16'h00d9,-16'h0513,16'h0126,16'h015a,16'h0141,16'h013a,16'h0006,-16'h0043,16'h000f,-16'h004b,-16'h012e,-16'h00bc,16'h0001,-16'h031e,16'h0088,-16'h009d,-16'h0219,-16'h0183,-16'h00de,-16'h0327,16'h014b,-16'h00bf,-16'h0351,-16'h018c,16'h0157,16'h00b9,-16'h037b,16'h0142,16'h003a,-16'h0081,16'h00ed,16'h0003,16'h00cf,-16'h003a,-16'h0011,16'h0188,16'h022d,16'h00f0,16'h0010,16'h0098,-16'h001d,16'h007c,16'h0102,-16'h0064,-16'h00ba,16'h0022,16'h009a,-16'h0009,16'h00f1,16'h0173,16'h0016,-16'h0083,-16'h051f,16'h0169,16'h0073,-16'h0160,16'h0031,16'h0023,-16'h003c,-16'h00a5,16'h00b3,-16'h01d2,-16'h00d2,-16'h00b8,16'h005e,-16'h0624,16'h015b,16'h0171,16'h018a,16'h01a7,16'h001a,-16'h0025,-16'h007c,-16'h009b,-16'h0117,-16'h00ce,-16'h0042,-16'h02b2,-16'h0006,-16'h0255,-16'h02f1,-16'h014e,-16'h0114,-16'h01d1,16'h0112,-16'h0064,-16'h076e,-16'h00bb,-16'h000f,16'h00f1,-16'h0391,16'h0141,16'h011d,-16'h0048,-16'h0024,-16'h0014,16'h0096,-16'h00ae,-16'h007b,16'h021c,16'h0279,16'h012c,-16'h0123,16'h00e9,16'h0016,16'h00b1,16'h0134,-16'h00a8,-16'h004f,16'h0040,16'h0028,-16'h005a,16'h0138,16'h00ba,16'h0045,-16'h005d,-16'h02f8,16'h004f,16'h00ac,-16'h01af,16'h003e,16'h0081,16'h0022,-16'h0101,16'h00ca,-16'h0231,-16'h00df,-16'h00e3,-16'h0028,-16'h04f3,16'h009c,16'h013f,16'h018c,16'h00d2,16'h0079,16'h0025,-16'h0057,-16'h0059,-16'h0122,-16'h008d,-16'h005f,-16'h016f,-16'h0216,-16'h027a,-16'h030c,-16'h0067,-16'h0103,-16'h0079,16'h00ed,-16'h003e,-16'h06a8,-16'h00b3,-16'h00bb,16'h013e,-16'h0298,16'h00d4,16'h0080,-16'h0072,-16'h009a,16'h0055,16'h00ec,16'h000b,16'h0021,16'h01a4,16'h02bc,16'h00e3,-16'h00f4,16'h004d,-16'h0078,16'h002c,16'h0105,-16'h0022,16'h0037,-16'h0081,16'h0045,-16'h003b,16'h0082,16'h005f,16'h004c,-16'h004b,-16'h0105,-16'h011b,16'h00c5,-16'h008d,16'h0130,16'h0028,-16'h0077,-16'h00c2,16'h008c,-16'h024c,-16'h0077,-16'h00d5,-16'h012d,-16'h03ae,-16'h0012,16'h00ef,16'h013c,16'h0118,16'h00cf,16'h00a0,-16'h0173,-16'h0054,-16'h0159,-16'h0083,16'h0071,-16'h0095,-16'h029e,-16'h0250,-16'h0280,-16'h005d,-16'h00e7,16'h00b4,16'h012c,16'h0000,-16'h0463,-16'h008a,-16'h0208,16'h0171,-16'h0184,16'h0045,16'h008a,16'h009c,-16'h0064,16'h0094,16'h000d,16'h00cf,16'h007a,16'h00e0,16'h02a5,-16'h00b4,-16'h01d9,-16'h005e,-16'h00af,-16'h0055,16'h00a5,16'h0023,16'h0017,-16'h000c,16'h000e,-16'h00a7,16'h0046,16'h010a,16'h0005,-16'h0051,-16'h007f,-16'h030b,16'h018c,-16'h00db,16'h0198,16'h000c,16'h00ec,16'h00b1,-16'h000f,-16'h004b,16'h0071,16'h0131,16'h00ba,16'h00fd,-16'h00d8,16'h0298,-16'h0013,16'h01c0,16'h012a,-16'h003c,16'h0039,-16'h00d9,-16'h0052,-16'h0013,-16'h0042,-16'h00d4,-16'h0045,16'h01b3,16'h0082,-16'h001c,-16'h023d,-16'h00f5,-16'h003f,-16'h01d1,16'h00b8,16'h02a1,16'h0089,16'h00b8,16'h0080,-16'h00ba,-16'h00aa,16'h006b,-16'h0002,-16'h005b,16'h023a,16'h0003,16'h0088,16'h0153,16'h0090,16'h00cd,-16'h00b0,16'h001b,16'h0005,16'h010f,-16'h00ac,16'h0023,-16'h0025,-16'h015f,-16'h0023,-16'h0209,16'h00ab,-16'h0020,-16'h0068,16'h0019,-16'h00d9,-16'h0170,-16'h0108,-16'h0058,16'h014f,-16'h0023,16'h00da,16'h0132,16'h0024,-16'h0081,16'h005d,16'h00b6,16'h0008,16'h0078,-16'h011d,16'h0118,-16'h00c0,16'h01de,16'h0196,-16'h0035,16'h0053,-16'h00de,16'h0043,16'h00d4,-16'h008e,16'h0046,-16'h0059,16'h005b,16'h00e8,-16'h0100,-16'h0323,-16'h014e,-16'h0046,-16'h0263,16'h00e8,16'h0240,16'h0074,16'h012d,16'h00b3,-16'h00e0,-16'h00e0,-16'h0017,16'h0062,-16'h0051,16'h022f,16'h00d2,16'h004a,16'h00b5,16'h014c,16'h0122,-16'h0035,16'h007e,16'h0011,16'h00d0,-16'h011e,-16'h003d,-16'h0047,-16'h004f,16'h00c1,-16'h01e2,16'h019c,16'h0018,-16'h0017,16'h00a8,-16'h0098,-16'h02e1,-16'h00b7,16'h0017,16'h0136,16'h004f,16'h01a6,16'h017a,16'h00c2,-16'h0037,-16'h0071,16'h008d,16'h000b,16'h0042,-16'h00e4,16'h011f,-16'h00ec,16'h0167,16'h0098,-16'h0010,16'h003d,-16'h0030,16'h00c8,16'h016a,-16'h00c6,16'h000c,-16'h017f,-16'h00d6,16'h0167,-16'h01af,-16'h0437,-16'h0067,-16'h0071,-16'h0284,16'h0059,16'h0165,16'h0067,16'h0100,16'h0061,16'h004b,-16'h00d2,16'h0004,16'h0032,16'h005b,16'h0191,16'h00d2,16'h0002,16'h0020,16'h013a,16'h00c9,-16'h006a,16'h0031,-16'h0021,16'h00a8,16'h0023,-16'h0008,16'h005e,-16'h00ce,16'h0088,-16'h0141,16'h01fd,-16'h007c,16'h0045,16'h003d,16'h003a,-16'h03e8,-16'h00ed,16'h0091,16'h007f,16'h0029,16'h01df,16'h00bd,16'h0146,-16'h0067,-16'h004c,16'h003a,16'h0056,16'h003c,-16'h00a2,16'h0031,-16'h02a2,16'h00eb,-16'h0123,-16'h004e,-16'h007f,16'h0071,16'h00be,16'h0171,-16'h00c9,16'h006a,-16'h015d,-16'h0059,16'h017c,-16'h01d2,-16'h0407,-16'h009a,16'h0007,-16'h02dd,-16'h0009,16'h0134,-16'h0036,16'h0065,-16'h005e,16'h013a,-16'h0050,-16'h0037,-16'h002b,16'h0163,16'h013a,16'h00a6,-16'h000c,16'h005b,16'h012f,16'h0118,-16'h0089,-16'h007e,-16'h00b0,16'h00a7,-16'h0052,16'h00cc,16'h0057,-16'h00f7,16'h012d,16'h003a,16'h0180,-16'h0137,-16'h004a,-16'h000d,16'h011d,-16'h03dd,-16'h0161,16'h0050,16'h0100,16'h0019,16'h0193,16'h0039,16'h018a,-16'h0074,-16'h0103,16'h0068,16'h0125,16'h001d,-16'h0113,16'h008b,-16'h0427,16'h0111,-16'h01a2,16'h0083,-16'h004a,16'h0016,16'h0109,16'h01cf,-16'h0028,16'h00bc,-16'h01ce,16'h003e,16'h01e0,-16'h0128,-16'h03b1,-16'h001f,-16'h0028,-16'h014f,16'h0029,16'h0174,16'h004f,16'h0003,-16'h00c6,16'h0224,-16'h0002,16'h0059,-16'h00b3,16'h0139,16'h0076,16'h0053,-16'h0067,16'h004b,16'h014d,16'h017b,-16'h00e3,-16'h0016,16'h002a,16'h0068,16'h0064,16'h0183,16'h0055,-16'h010d,16'h00dd,16'h0114,16'h014f,-16'h0034,-16'h006d,-16'h00cb,16'h016c,-16'h0489,-16'h00e4,16'h002d,16'h0113,16'h0042,16'h0134,16'h0079,16'h01f9,-16'h0027,-16'h00f9,-16'h0032,16'h01b7,16'h003f,-16'h00dc,16'h00f6,-16'h0531,16'h01b3,-16'h015b,16'h0066,-16'h0057,16'h000d,16'h00bf,16'h01ff,-16'h0010,16'h00ff,-16'h0157,-16'h0004,16'h02ac,16'h002d,-16'h0281,16'h0009,16'h006f,-16'h0014,16'h000e,16'h00f0,-16'h0099,-16'h0053,-16'h01a1,16'h0218,16'h007e,-16'h000d,-16'h0083,16'h0102,-16'h0039,-16'h004a,16'h0027,-16'h0052,16'h01fb,16'h0105,-16'h013c,16'h008e,16'h0076,-16'h0038,16'h006f,16'h01a1,16'h004a,-16'h00ff,16'h00eb,16'h010c,16'h00ad,-16'h002d,-16'h00fc,-16'h00ea,16'h0182,-16'h047b,-16'h0084,16'h00b1,16'h00ae,16'h0067,16'h0105,16'h006f,16'h0234,-16'h0043,-16'h0084,16'h0033,16'h01e9,16'h0049,-16'h00ca,16'h00bd,-16'h034c,16'h0173,-16'h0093,16'h004c,-16'h00c2,-16'h006d,16'h00ba,16'h0214,16'h0001,16'h0153,16'h000d,16'h003a,16'h0350,16'h0251,-16'h0267,16'h0050,16'h0080,-16'h0030,16'h0075,16'h015e,-16'h009f,16'h0045,-16'h0101,16'h01ff,-16'h00dc,-16'h0055,-16'h002a,16'h0096,-16'h0045,-16'h00c5,-16'h0057,-16'h0020,16'h019c,16'h00f4,-16'h009a,16'h00e5,16'h0072,16'h0001,16'h0023,16'h01b4,16'h0010,-16'h00f2,16'h00be,16'h00f2,-16'h0074,16'h000f,-16'h0131,-16'h00bd,16'h01f4,-16'h0441,-16'h0063,16'h006d,16'h0131,16'h0033,16'h008a,16'h0099,16'h0168,-16'h0010,-16'h0071,16'h0080,16'h020b,16'h0096,-16'h00f1,16'h0122,-16'h02a8,16'h01d2,16'h0098,16'h008d,-16'h0002,16'h0005,16'h007b,16'h0258,-16'h003c,-16'h0065,16'h0085,16'h0080,16'h0257,16'h0299,-16'h027f,16'h00bf,16'h00d5,-16'h01f8,16'h005e,16'h01a1,16'h0042,16'h0091,16'h0060,16'h005d,-16'h0113,-16'h004a,16'h0169,16'h0032,-16'h00bb,-16'h00d4,-16'h01b4,16'h0095,16'h01a5,16'h0117,-16'h005b,16'h015e,16'h0056,16'h00aa,-16'h005f,16'h022c,16'h0013,-16'h00d8,16'h00ec,16'h019d,-16'h0154,16'h008b,-16'h00c6,16'h00b9,16'h0196,-16'h0424,-16'h0060,-16'h0021,16'h009e,16'h0045,16'h002c,16'h0030,16'h01f4,-16'h0040,-16'h00ba,16'h00db,16'h017d,16'h00d6,-16'h00a7,16'h01bc,-16'h01b0,16'h01cf,16'h0060,16'h0116,-16'h002f,-16'h0088,16'h009a,16'h01ff,16'h0022,-16'h004f,16'h0136,16'h015b,16'h020b,16'h0152,-16'h0203,16'h009e,16'h0114,-16'h037a,16'h00a0,16'h0065,16'h019a,16'h00e7,16'h0074,-16'h0132,-16'h0072,-16'h002e,16'h01ec,16'h00ac,-16'h0113,16'h007e,-16'h0255,16'h00e3,16'h01a8,16'h018c,16'h0024,16'h00dc,16'h0084,16'h00d8,-16'h00cc,16'h0268,-16'h0092,-16'h00a4,16'h00dd,16'h0201,-16'h01f0,16'h0107,-16'h0085,16'h0129,16'h0200,-16'h0334,-16'h0039,-16'h002e,16'h0102,16'h002d,-16'h006d,16'h0051,16'h017b,-16'h0074,-16'h000b,16'h0080,16'h01c3,16'h00e2,-16'h0090,16'h00fe,-16'h0075,16'h0166,16'h0017,16'h01c2,-16'h000e,-16'h00c8,16'h00db,16'h01bf,16'h0089,16'h004d,16'h01e8,16'h00c4,16'h0105,16'h00e9,-16'h01e6,16'h007f,16'h0178,-16'h033b,16'h0088,-16'h009b,16'h0209,16'h0114,16'h0089,-16'h012c,16'h0107,-16'h0050,16'h000e,16'h003d,-16'h00b7,16'h01b5,-16'h0181,16'h00a0,16'h021a,16'h0185,16'h009c,16'h0094,16'h0060,16'h0061,-16'h0197,16'h025f,-16'h004b,-16'h00db,-16'h0073,16'h012a,-16'h00cb,16'h00b8,16'h0082,16'h00e9,16'h0254,-16'h01fb,-16'h0051,16'h0004,16'h0102,16'h006b,-16'h0028,16'h0098,16'h01bb,-16'h009e,-16'h0069,16'h00bb,16'h0184,16'h009d,-16'h0018,16'h001d,16'h0152,16'h0168,16'h0000,16'h012f,-16'h0029,-16'h0103,16'h011c,16'h01bf,16'h00be,-16'h001f,16'h0199,16'h00e6,16'h011b,-16'h010e,-16'h01b4,16'h0069,16'h0163,-16'h00df,16'h0081,-16'h014b,16'h0259,16'h00c1,16'h00a7,-16'h0044,16'h015d,16'h0003,-16'h01e1,-16'h0027,-16'h00d0,16'h0101,16'h00a1,16'h005f,16'h01d9,16'h010c,16'h00ae,16'h0007,16'h002f,16'h0080,-16'h021f,16'h0242,-16'h0004,-16'h0087,-16'h0028,16'h0114,16'h0092,16'h0135,16'h0144,16'h00b9,16'h025e,-16'h01b3,-16'h0026,16'h007c,16'h008b,-16'h0001,16'h001b,16'h0078,16'h01b0,16'h0013,-16'h005a,16'h00cf,16'h00fc,16'h0067,-16'h0028,16'h012b,16'h0264,16'h0134,-16'h00de,16'h004c,-16'h0068,-16'h0124,16'h0127,16'h015b,16'h00af,16'h005f,16'h00f1,16'h0024,16'h0154,-16'h020e,-16'h014e,-16'h003d,16'h00d8,16'h0082,16'h0083,-16'h0152,16'h017e,16'h0096,16'h00f1,16'h0068,16'h005f,-16'h004f,-16'h0229,16'h0057,-16'h0010,16'h00ad,16'h00fa,16'h007e,16'h015c,16'h011c,16'h00fd,16'h0077,-16'h0012,16'h0037,-16'h00fd,16'h01ef,16'h0099,-16'h0125,-16'h00b5,16'h007f,16'h0134,16'h0138,16'h00d3,16'h00c5,16'h0203,-16'h0198,16'h0024,16'h0069,16'h00a0,16'h0034,16'h009b,-16'h0043,16'h01f1,16'h0070,-16'h00e4,16'h0098,16'h0120,-16'h006d,16'h0051,16'h0050,16'h0209,16'h009e,-16'h00b2,-16'h0013,-16'h0088,-16'h00b1,16'h0140,16'h012d,-16'h000f,16'h00b8,16'h00aa,-16'h00cf,16'h009e,-16'h02a5,-16'h0201,-16'h00e6,16'h0149,16'h0052,-16'h006e,-16'h003f,16'h0032,16'h006d,16'h0161,16'h01d8,-16'h004e,-16'h0051,-16'h019d,16'h0039,16'h0035,16'h0035,16'h00dc,16'h0016,16'h0116,16'h00c8,16'h00e9,16'h008c,16'h0019,16'h00ad,-16'h007b,16'h01a3,16'h00a4,-16'h00c2,-16'h010a,16'h00cf,16'h0213,16'h00ff,16'h0113,16'h0115,16'h01fb,-16'h007b,16'h00a4,16'h0081,16'h00e1,16'h0010,16'h0066,16'h0005,16'h01bf,16'h0026,-16'h006b,16'h00da,16'h005b,-16'h00c4,16'h0036,-16'h006c,16'h0191,16'h00e0,-16'h0060,-16'h007b,-16'h0070,-16'h00e6,16'h014e,16'h006d,16'h004b,16'h0085,16'h003b,-16'h00f8,16'h010c,-16'h0285,-16'h017c,16'h00fa,16'h00ee,16'h000b,-16'h00ff,16'h00bf,-16'h0112,16'h007f,16'h00ee,16'h01e1,-16'h00c4,-16'h0011,16'h0111,16'h0016,-16'h0018,16'h000e,16'h00cd,16'h0101,16'h00bd,16'h0134,16'h0124,16'h0093,-16'h0016,16'h0089,-16'h0049,16'h00f4,16'h0010,-16'h00ab,-16'h002c,16'h006f,16'h0227,16'h011d,16'h0197,16'h00e4,16'h0201,16'h003e,16'h00bb,16'h0019,16'h0096,16'h0089,16'h00c3,16'h0046,16'h010f,16'h0051,-16'h0064,16'h0046,-16'h0020,-16'h0003,16'h006b,16'h004d,16'h01be,16'h00f8,16'h0019,-16'h0021,-16'h005e,-16'h013d,16'h0135,16'h007a,16'h00af,16'h0098,16'h007e,16'h000d,16'h01b8,-16'h022c,-16'h0045,16'h01ea,16'h0107,-16'h001d,-16'h012e,16'h014b,-16'h02c8,16'h00b1,16'h005a,16'h01ae,-16'h006e,-16'h007c,16'h012a,16'h007d,-16'h0075,16'h0128,-16'h0004,16'h017b,16'h0089,16'h00a6,16'h0085,16'h00ed,16'h002e,16'h004f,-16'h0035,16'h0129,-16'h004c,-16'h010c,-16'h00ec,16'h00b0,-16'h0070,16'h00ce,16'h01e0,16'h0063,16'h021e,16'h00ee,16'h00e8,-16'h0033,16'h0094,16'h0065,16'h0164,16'h00e6,16'h0112,16'h0020,-16'h0097,16'h0014,-16'h002d,16'h001e,-16'h0029,16'h00f4,16'h01ad,16'h009c,16'h0030,16'h0032,-16'h0043,-16'h0156,16'h0184,16'h0071,16'h0016,16'h00a6,-16'h0032,16'h001a,16'h01d0,-16'h0043,16'h0068,16'h018b,16'h013e,-16'h00ba,-16'h0190,16'h00fb,-16'h0227,16'h00a2,16'h008f,16'h00ad,16'h003f,16'h0008,16'h00b0,16'h0112,-16'h00b7,16'h00b6,16'h00b5,16'h013b,16'h00e9,16'h0118,16'h00ba,16'h00db,16'h0066,16'h0048,-16'h0092,16'h0191,-16'h0009,-16'h005e,-16'h00e0,16'h00cc,-16'h0185,16'h0126,16'h01ac,16'h00b7,16'h024c,16'h014b,16'h0118,16'h002e,16'h009f,16'h00ae,16'h015d,16'h0078,16'h0093,16'h005e,-16'h0105,16'h0028,-16'h000c,-16'h003a,16'h0003,16'h00fc,16'h0142,16'h00e4,16'h001d,16'h004a,16'h0014,-16'h0118,16'h0202,16'h004e,-16'h001e,16'h0049,-16'h003a,16'h0049,16'h006d,16'h007b,16'h0000,16'h0206,16'h0119,-16'h0138,-16'h00f5,16'h002c,-16'h021f,16'h0090,-16'h003a,16'h005d,16'h0048,16'h005d,16'h00bb,16'h0034,-16'h0182,16'h0027,16'h005b,16'h012b,16'h007a,16'h00f2,16'h002b,16'h0039,16'h0037,16'h00b5,16'h0099,16'h01ce,16'h0009,-16'h0021,-16'h001f,16'h0049,-16'h0239,16'h0126,16'h01c9,16'h006d,16'h01b0,16'h00bb,16'h0128,-16'h00cd,16'h00fa,16'h001d,16'h013a,16'h00a9,16'h011c,16'h0027,16'h004d,16'h0106,-16'h0007,16'h000c,16'h0036,16'h0012,16'h00e1,16'h00bd,16'h003e,16'h00bd,-16'h0015,-16'h00fa,16'h026c,16'h008a,-16'h0016,16'h00c2,-16'h00bd,16'h0042,-16'h001a,16'h00f4,-16'h0087,16'h020d,16'h014d,-16'h00f4,16'h00e8,-16'h00cb,-16'h025b,16'h0019,-16'h0078,-16'h0024,16'h0094,16'h0088,-16'h0059,-16'h003f,-16'h0173,16'h0010,16'h0074,16'h0119,16'h0080,16'h00c6,16'h0025,-16'h0058,16'h0013,16'h0104,16'h0084,16'h01e1,16'h0021,-16'h0063,16'h0012,16'h003a,-16'h0135,16'h01bc,16'h015c,16'h0045,16'h01c1,16'h0106,16'h0136,-16'h017c,16'h00f8,16'h007c,16'h002f,16'h0063,16'h00ea,16'h0009,16'h00eb,16'h00a3,16'h0083,-16'h0030,16'h010e,-16'h000c,16'h0055,16'h00a3,-16'h0010,16'h0028,-16'h003a,-16'h0094,16'h0207,16'h00b1,-16'h005e,16'h00a3,-16'h00b9,16'h006a,-16'h00fc,16'h012f,16'h0012,16'h015c,16'h01e0,-16'h0090,16'h0182,-16'h00de,-16'h00e6,16'h0024,16'h00a7,-16'h0094,16'h006c,16'h00a9,-16'h0098,-16'h0037,-16'h00f8,16'h0063,16'h01a8,16'h013b,16'h00b0,16'h00e2,16'h008e,-16'h0004,16'h0071,16'h002d,16'h0050,16'h018e,-16'h0062,-16'h011b,-16'h003b,16'h003a,16'h006c,16'h013e,16'h011a,16'h0037,16'h01f9,16'h0088,16'h0105,-16'h0143,16'h0129,16'h0040,16'h0085,-16'h0017,16'h00f7,16'h0049,16'h0108,-16'h0023,16'h00ee,-16'h00b5,16'h0037,16'h0050,16'h000a,16'h008d,-16'h002f,16'h0046,16'h00c3,-16'h005d,16'h016f,16'h00b5,-16'h0012,16'h007b,-16'h0082,16'h00a4,-16'h00a5,16'h0146,-16'h0084,16'h00cb,16'h01b3,-16'h0082,16'h01ad,-16'h00b7,-16'h0075,16'h0012,16'h00c6,-16'h005f,-16'h0054,16'h0035,-16'h002d,-16'h0004,-16'h006e,16'h0059,16'h00d4,16'h00d3,16'h011b,16'h00ee,16'h00ba,-16'h0023,16'h0070,16'h0028,16'h0005,16'h01c1,-16'h0007,-16'h00cc,-16'h001b,16'h000d,16'h00c6,16'h00e7,16'h00fb,-16'h0013,16'h024e,-16'h000a,16'h0087,-16'h017f,16'h0089,16'h0025,-16'h001c,16'h005c,16'h010b,16'h00d6,16'h0115,-16'h0081,16'h00a3,-16'h0050,16'h0018,16'h0065,-16'h00aa,16'h00c0,-16'h00a5,16'h0078,16'h009b,-16'h00cf,16'h0139,16'h0053,-16'h0055,16'h0178,16'h0045,16'h00c2,-16'h00b2,16'h00ea,-16'h001f,-16'h02c7,16'h0187,-16'h012a,16'h01f1,-16'h00c5,16'h009c,16'h010c,16'h015e,-16'h0053,-16'h00c8,16'h0054,-16'h007f,-16'h0059,-16'h0010,16'h008e,16'h00cf,16'h00dd,16'h0070,16'h011c,-16'h0001,16'h004a,-16'h0041,16'h00a0,-16'h0009,16'h00fb,-16'h00bf,-16'h005f,16'h0037,-16'h0097,16'h004a,16'h0100,16'h00c1,-16'h009a,16'h0257,16'h0036,16'h0018,-16'h0076,16'h014e,-16'h0089,-16'h0072,16'h008d,16'h00cf,16'h008b,16'h0148,-16'h009a,16'h0088,-16'h0166,-16'h0024,16'h0101,-16'h013e,16'h0131,16'h0047,16'h006e,16'h0060,-16'h00a3,16'h0164,16'h0017,-16'h0022,16'h00eb,16'h0093,16'h0139,-16'h00fb,16'h00d8,-16'h014c,-16'h08e9,16'h00cd,-16'h00de,16'h0188,-16'h0036,16'h00c2,16'h005b,16'h00a5,16'h009b,-16'h00bd,-16'h0026,-16'h004e,-16'h003a,16'h00de,16'h00df,16'h00cd,16'h013a,16'h0097,16'h00af,-16'h00e2,-16'h0030,16'h0036,16'h00ff,16'h003a,16'h0131,-16'h008a,-16'h00c4,16'h0021,-16'h00a1,16'h00b9,16'h00d3,16'h0034,-16'h0055,16'h0151,16'h0070,16'h0045,16'h0024,16'h0118,-16'h009a,-16'h00ee,16'h0008,16'h008b,16'h009b,-16'h0013,-16'h00cd,16'h0060,-16'h03de,16'h0084,16'h00eb,16'h0067,16'h00f9,-16'h0016,-16'h002c,16'h0007,-16'h00b0,16'h0097,-16'h0017,16'h0006,-16'h00e6,16'h00ee,16'h00de,-16'h012a,16'h0098,-16'h01cf,-16'h0a00,16'h015b,-16'h00c7,16'h016a,-16'h002d,16'h0118,16'h0026,-16'h0001,16'h0105,-16'h0046,-16'h0015,-16'h0008,-16'h0051,16'h00ed,16'h008c,16'h0151,16'h01b6,16'h012b,16'h0048,-16'h00da,16'h001e,16'h0043,16'h0044,16'h002a,16'h0169,-16'h00b1,-16'h010b,-16'h0014,-16'h018a,16'h00e8,16'h0144,16'h0008,16'h0001,-16'h0236,16'h005e,16'h00c1,16'h0009,16'h00a8,-16'h00ae,-16'h0086,-16'h007b,16'h00e1,-16'h0005,-16'h0077,-16'h0107,16'h00e2,-16'h05cf,16'h00c8,16'h0129,16'h0105,16'h00cb,16'h0027,-16'h0001,16'h0017,-16'h00ae,16'h00e7,-16'h0043,-16'h001b,-16'h0319,16'h0136,-16'h0056,-16'h01a6,-16'h00c0,-16'h014f,-16'h056e,16'h00db,-16'h006a,16'h0096,-16'h00ea,16'h0150,16'h0048,-16'h016a,16'h01a0,-16'h0028,-16'h0081,16'h0115,-16'h0053,16'h009c,16'h00bb,16'h005a,16'h00f9,16'h0130,16'h008d,-16'h004c,16'h00c3,-16'h0002,16'h0033,-16'h0053,16'h014c,-16'h00af,16'h0006,16'h002a,-16'h00fe,16'h0143,16'h012f,-16'h0019,16'h0055,-16'h06ae,16'h00ba,16'h0055,-16'h0089,16'h0011,-16'h005a,-16'h00d4,-16'h00bc,16'h00f5,16'h0025,-16'h011e,-16'h010a,16'h0129,-16'h06e5,16'h0147,16'h01a9,16'h01a1,16'h00d4,16'h00ae,16'h0047,16'h0039,-16'h0114,16'h00b0,16'h002e,16'h001b,-16'h02c8,16'h00ce,-16'h01ff,-16'h01fa,-16'h01bc,-16'h00a4,-16'h036e,16'h012c,-16'h0099,-16'h036b,-16'h0131,16'h0094,16'h0086,-16'h027c,16'h014a,16'h00a2,-16'h0083,16'h00bc,-16'h0048,16'h00ad,-16'h0013,-16'h0012,16'h0187,16'h020e,16'h00a5,-16'h00c9,16'h0104,16'h0052,16'h0080,16'h00b5,-16'h0018,-16'h0007,16'h005c,-16'h0071,16'h001c,16'h00df,16'h012d,16'h0001,16'h0001,-16'h06c5,16'h014e,16'h006f,-16'h0109,16'h001f,-16'h0008,16'h0009,-16'h011d,16'h009f,-16'h00d6,-16'h00ac,-16'h00e1,16'h00a8,-16'h0546,16'h015c,16'h01a1,16'h01b3,16'h009e,16'h0010,-16'h003c,-16'h006b,-16'h007c,16'h005a,-16'h0024,-16'h003c,-16'h0227,-16'h00bd,-16'h02ae,-16'h023d,-16'h00bb,-16'h0189,-16'h019b,16'h016f,-16'h007b,-16'h0739,-16'h00c2,-16'h0067,16'h0070,-16'h01fc,16'h0107,16'h00ec,16'h0055,16'h0039,-16'h0025,16'h008a,16'h002b,-16'h003f,16'h023a,16'h0220,16'h0084,-16'h00e7,16'h00b1,-16'h000a,16'h0086,16'h0125,16'h0001,-16'h0067,-16'h0020,16'h005c,16'h0021,16'h0070,16'h00df,16'h0097,-16'h0009,-16'h03af,-16'h003c,16'h00ac,-16'h01a0,16'h012c,16'h001f,16'h005f,-16'h0125,16'h0117,-16'h0227,-16'h0035,-16'h00d8,-16'h006b,-16'h0453,16'h012f,16'h0171,16'h0168,16'h00b9,16'h0096,16'h000c,-16'h010b,-16'h0023,-16'h0002,-16'h000b,-16'h0015,-16'h00fa,-16'h01dd,-16'h030c,-16'h02a7,16'h0012,-16'h0111,-16'h0039,16'h012e,-16'h001c,-16'h065a,-16'h0002,-16'h01be,16'h005d,-16'h015d,16'h006d,16'h00c4,16'h0025,16'h004f,16'h003d,16'h0035,16'h0016,-16'h0053,16'h025f,16'h021d,16'h0075,-16'h019a,16'h003b,-16'h0057,16'h0017,16'h0115,-16'h0032,16'h0062,16'h0051,16'h00aa,16'h000e,16'h0040,16'h009b,16'h00e3,16'h00a4,-16'h01ad,-16'h0113,16'h006e,-16'h0063,16'h00e9,-16'h001f,16'h0067,-16'h00fb,16'h008b,-16'h02bb,-16'h0016,-16'h0130,-16'h012e,-16'h03a1,16'h0000,16'h00c9,16'h012c,16'h008e,16'h00de,16'h00c0,-16'h0186,-16'h003a,16'h0022,-16'h0038,16'h0008,-16'h001e,-16'h0229,-16'h0212,-16'h01d2,-16'h0078,-16'h00d0,16'h00b8,16'h01cc,16'h0080,-16'h042c,16'h0010,-16'h0252,16'h018b,-16'h00c3,16'h0011,16'h003f,16'h007c,16'h0027,16'h00b2,16'h005b,16'h0095,16'h009f,16'h01c6,16'h02eb,-16'h00c2,-16'h0208,-16'h00a3,-16'h00c8,-16'h005d,16'h014c,16'h004f,16'h005d,-16'h0004,16'h0080,-16'h009b,16'h0047,16'h00db,16'h000b,16'h0047,-16'h0121,-16'h0208,16'h00d0,-16'h002e,16'h016f,16'h0024,16'h015b,16'h012b,-16'h0024,16'h000d,16'h00cf,16'h0111,16'h00c0,16'h011a,-16'h00b0,16'h02da,-16'h00d8,16'h01b9,16'h00c8,-16'h0001,16'h0066,-16'h0083,-16'h00a2,16'h0000,-16'h001b,-16'h00da,16'h0039,16'h023f,-16'h0007,16'h0001,-16'h0274,-16'h01a3,16'h000a,-16'h0101,16'h00a2,16'h0335,16'h018d,16'h00bc,16'h00ec,-16'h0101,-16'h00d7,-16'h000e,-16'h0041,-16'h0068,16'h029e,-16'h007d,16'h0066,16'h0186,16'h00ad,16'h000b,-16'h0012,16'h003b,16'h0019,16'h0109,-16'h0128,16'h004a,-16'h0021,-16'h00bb,16'h00d8,-16'h01d2,16'h0094,16'h0039,-16'h0113,-16'h0006,-16'h0091,-16'h00a5,-16'h00fc,16'h00c6,16'h0116,16'h000e,16'h0161,16'h0192,16'h0035,-16'h00e7,16'h00b0,16'h008d,16'h0071,16'h00d0,16'h0026,16'h0210,-16'h0122,16'h01e6,16'h00cd,16'h004f,16'h004c,-16'h00b5,16'h0019,16'h007a,-16'h00a2,-16'h003e,-16'h007b,16'h002e,16'h0127,-16'h00d4,-16'h032f,-16'h00ae,-16'h00ac,-16'h0187,16'h0076,16'h01b9,16'h00ff,16'h0109,16'h0106,-16'h0105,-16'h00bc,-16'h0085,-16'h0005,16'h001a,16'h022f,16'h003e,16'h0023,16'h0147,16'h014a,16'h0073,16'h0009,16'h0096,-16'h004e,16'h00ad,-16'h00e8,-16'h0015,-16'h002a,-16'h0042,16'h00a0,-16'h0153,16'h0117,-16'h0050,-16'h001a,16'h0034,-16'h00a4,-16'h01d2,-16'h0136,16'h0059,16'h012f,16'h0082,16'h0188,16'h01c8,-16'h0052,-16'h00f4,16'h0052,16'h00ac,-16'h0009,16'h0057,16'h008e,16'h0164,-16'h0199,16'h01aa,16'h0021,16'h0056,16'h002b,16'h0001,16'h009a,16'h0148,-16'h0088,-16'h000a,-16'h012f,-16'h00bc,16'h0155,-16'h0144,-16'h03fc,-16'h0070,-16'h00d0,-16'h0245,16'h0031,16'h0164,16'h005c,16'h00b5,16'h0070,-16'h0006,-16'h0079,-16'h0096,-16'h0057,16'h00b2,16'h017c,16'h00bf,-16'h0033,16'h00ba,16'h0169,16'h00ed,16'h004d,16'h0060,16'h0036,16'h0050,-16'h00b3,16'h0014,-16'h0014,-16'h0099,16'h00f6,-16'h001b,16'h0185,-16'h0049,16'h0004,-16'h0074,-16'h0066,-16'h01dd,-16'h0198,-16'h000d,16'h00af,16'h0036,16'h0194,16'h0132,-16'h0044,-16'h007b,-16'h000d,16'h0015,-16'h0066,16'h0064,16'h0005,16'h002d,-16'h029d,16'h013c,-16'h0054,16'h002d,-16'h0007,16'h001b,16'h00b9,16'h016f,-16'h0109,16'h0003,-16'h01d8,-16'h0068,16'h0162,-16'h010b,-16'h0421,-16'h007c,-16'h00b4,-16'h0168,-16'h006e,16'h0104,-16'h0079,16'h0072,-16'h0091,16'h0100,-16'h000c,-16'h0132,-16'h0027,16'h00e2,16'h0187,16'h0095,16'h0004,16'h004c,16'h019b,16'h00e9,16'h001c,16'h0083,16'h0004,16'h00e1,-16'h0021,16'h00de,16'h0087,-16'h0120,16'h00ff,16'h015f,16'h015c,-16'h010e,-16'h0064,-16'h0048,16'h00a1,-16'h01f4,-16'h01f7,-16'h005b,16'h00a1,16'h001f,16'h017d,16'h00b7,-16'h0053,-16'h002b,-16'h0061,16'h00c1,16'h0148,16'h003c,16'h0042,16'h000b,-16'h0374,16'h0129,-16'h00ef,16'h003a,-16'h0063,16'h0009,16'h0092,16'h01cc,-16'h00d1,16'h0124,-16'h0282,16'h0011,16'h0224,-16'h0043,-16'h0360,16'h0051,-16'h0043,-16'h00e4,-16'h0032,16'h0183,16'h0000,16'h0038,-16'h024f,16'h0210,16'h00a8,-16'h00dc,-16'h0031,16'h00d0,16'h011e,16'h0009,16'h0053,16'h003e,16'h01ae,16'h00ba,-16'h0030,16'h005e,16'h005c,16'h00ac,-16'h0014,16'h0157,16'h0043,-16'h00c3,16'h00f5,16'h01a1,16'h0153,-16'h0089,-16'h007f,-16'h00cd,16'h00e5,-16'h01cc,-16'h01d2,16'h0029,16'h00f1,16'h0009,16'h0174,16'h015c,16'h0010,-16'h0016,16'h0020,16'h0074,16'h0149,-16'h0012,-16'h000d,16'h00c4,-16'h03fb,16'h00bd,-16'h00f6,16'h000b,-16'h0057,-16'h0098,16'h0061,16'h0248,-16'h0086,16'h00d6,-16'h023f,16'h003e,16'h02c7,16'h00dd,-16'h02a4,16'h00af,16'h0069,-16'h006d,16'h0028,16'h010a,-16'h0006,16'h00eb,-16'h01bc,16'h01ef,-16'h0039,-16'h007a,-16'h00b8,16'h0119,16'h000e,-16'h001a,16'h0001,-16'h00ae,16'h0200,16'h009d,-16'h0069,16'h0127,16'h00a3,16'h0063,-16'h0012,16'h0197,16'h0090,-16'h009e,16'h00c2,16'h01da,-16'h0042,-16'h004f,-16'h0151,-16'h00f6,16'h012f,-16'h0190,-16'h01f1,-16'h0028,16'h00f5,16'h003f,16'h011c,16'h00f0,16'h0018,16'h0010,16'h000d,16'h001f,16'h018c,16'h0016,-16'h0016,16'h0124,-16'h037d,16'h0147,-16'h0065,-16'h000f,-16'h000b,-16'h0086,16'h008a,16'h020b,-16'h0095,16'h00f2,-16'h005f,16'h0058,16'h0265,16'h020c,-16'h027d,16'h00c5,16'h003f,-16'h016b,16'h0055,16'h0181,16'h0075,16'h007b,-16'h0132,16'h01ca,-16'h016d,-16'h00bc,16'h0038,16'h0080,-16'h0086,-16'h0027,-16'h0072,-16'h0042,16'h0201,16'h00ed,-16'h0034,16'h012a,16'h00ff,16'h006e,-16'h0069,16'h0143,16'h0014,-16'h0039,16'h00f1,16'h01df,-16'h00c6,16'h0076,-16'h01aa,-16'h00f5,16'h018f,-16'h017f,-16'h016c,16'h0063,16'h0087,16'h0064,16'h00c6,16'h00d9,-16'h0024,-16'h001f,16'h00c8,16'h009a,16'h01ce,16'h0091,-16'h006d,16'h0177,-16'h01f5,16'h0197,-16'h0032,16'h0061,16'h003b,16'h0024,16'h0085,16'h020c,-16'h0023,-16'h0023,16'h005f,16'h0060,16'h0251,16'h0240,-16'h0264,16'h00d4,16'h0090,-16'h0253,16'h0082,16'h01e9,16'h015c,16'h00a6,16'h0078,16'h001e,-16'h0172,-16'h005a,16'h0171,16'h0020,-16'h003c,-16'h0044,-16'h0184,-16'h0055,16'h0187,16'h0119,-16'h004e,16'h005e,16'h00e7,16'h0077,-16'h005b,16'h01df,-16'h006a,-16'h00a8,16'h009f,16'h027c,-16'h00b7,16'h00e8,-16'h00f5,16'h005c,16'h018a,-16'h015a,-16'h01a1,-16'h005d,16'h00f1,-16'h002e,16'h0065,16'h0090,-16'h0087,-16'h004c,16'h0078,16'h0068,16'h0129,16'h008b,-16'h005c,16'h01de,-16'h006a,16'h0171,-16'h0016,16'h0108,-16'h0089,-16'h007d,16'h00b9,16'h024f,16'h0089,-16'h0024,16'h016f,16'h00c7,16'h01b6,16'h017e,-16'h01f8,16'h0094,16'h0086,-16'h03bb,16'h002e,16'h00cb,16'h0286,16'h00f2,16'h002d,-16'h00f1,-16'h0090,-16'h009e,16'h01d5,16'h0058,-16'h00cd,16'h0119,-16'h021d,-16'h001b,16'h0164,16'h0128,16'h00e7,16'h0045,16'h00fb,16'h00f0,-16'h013a,16'h021a,16'h0031,-16'h002a,16'h0000,16'h01ef,-16'h021f,16'h0116,-16'h00f2,16'h00a7,16'h0119,-16'h0025,-16'h0210,-16'h00ce,16'h0119,-16'h0062,16'h0052,16'h0091,-16'h0069,-16'h0003,16'h00b9,16'h005d,16'h00ce,16'h0037,-16'h0079,16'h0112,16'h00ab,16'h00f1,-16'h006c,16'h01cb,-16'h006c,-16'h001c,16'h0120,16'h012a,16'h00c4,-16'h0058,16'h01f1,16'h0153,16'h0155,16'h005f,-16'h0196,16'h0088,16'h00fe,-16'h036a,16'h0016,-16'h0190,16'h01f6,16'h00ce,16'h0085,-16'h00ca,16'h0178,-16'h0073,-16'h002d,-16'h0020,-16'h00b7,16'h0186,-16'h0159,-16'h0004,16'h020c,16'h019d,16'h0119,16'h00f7,16'h00a0,16'h00be,-16'h0133,16'h0257,16'h0044,16'h0015,-16'h013f,16'h00e0,-16'h0162,16'h009c,-16'h001d,16'h003c,16'h01cd,16'h004f,-16'h017f,-16'h008b,16'h00f5,-16'h0041,16'h00e3,16'h00da,16'h0062,16'h0021,16'h005c,16'h00c1,16'h0106,16'h004c,-16'h0057,16'h00dd,16'h01c8,16'h00e0,-16'h00ed,16'h018f,-16'h0079,-16'h0042,16'h00f3,16'h009a,16'h003c,-16'h0043,16'h01cc,16'h0103,16'h013f,-16'h0204,-16'h0102,16'h0001,16'h0111,-16'h0007,16'h00d2,-16'h0262,16'h0168,16'h00d4,16'h0048,-16'h003a,16'h0142,16'h0073,-16'h0264,16'h0029,-16'h0082,16'h01cf,-16'h0057,-16'h0012,16'h015f,16'h0129,16'h00ef,16'h0048,16'h00b0,16'h0024,-16'h0149,16'h024a,16'h0077,16'h0052,-16'h00fd,16'h000f,16'h0090,16'h00ed,16'h0099,-16'h0028,16'h017e,16'h0032,-16'h01b6,-16'h009d,16'h00c5,-16'h0017,16'h0083,16'h0070,16'h00d8,16'h00a7,-16'h000d,16'h00f6,16'h00c2,16'h0071,-16'h009f,16'h0099,16'h01b3,16'h011f,-16'h00be,16'h0089,-16'h0070,-16'h00a8,16'h00c8,16'h00dc,16'h0009,-16'h0064,16'h0170,-16'h0070,16'h00ff,-16'h020e,-16'h0152,-16'h0078,16'h0125,16'h0126,16'h0114,-16'h01cd,16'h00ac,16'h0105,16'h003b,16'h008d,16'h00d8,-16'h003d,-16'h02c5,-16'h000f,16'h0019,16'h010f,16'h00cd,16'h0001,16'h0101,16'h0137,16'h00e1,16'h006c,16'h00dc,-16'h0018,-16'h0109,16'h0219,16'h012f,-16'h00db,-16'h0149,16'h003e,16'h0128,16'h009c,16'h0069,16'h006d,16'h0143,16'h0030,-16'h01be,-16'h0137,16'h0111,-16'h0033,16'h008f,16'h00c4,16'h00ca,16'h00ea,-16'h0086,16'h0107,16'h00fb,16'h002f,-16'h00d2,16'h0028,16'h0124,16'h00bb,-16'h002a,-16'h0011,-16'h0036,-16'h000b,16'h011b,16'h0127,-16'h003c,16'h00e0,16'h0077,-16'h0107,16'h018c,-16'h0238,-16'h0136,-16'h00bb,16'h0167,16'h008f,16'h0026,-16'h00e6,-16'h00b6,16'h00ba,16'h00ef,16'h0157,-16'h0021,16'h005d,-16'h0193,16'h002f,16'h00c2,-16'h0008,16'h0011,16'h0094,16'h00a5,16'h00bc,16'h00e1,16'h0080,16'h0065,16'h001f,-16'h011b,16'h0209,16'h00fc,-16'h00e5,-16'h018f,16'h0019,16'h0228,16'h0114,16'h00a6,16'h0068,16'h011b,16'h0055,-16'h0124,-16'h0090,16'h0161,-16'h0050,16'h00ce,16'h009f,16'h0076,16'h008f,-16'h000d,16'h007b,16'h00e7,16'h0044,-16'h003d,-16'h0014,16'h0134,16'h00b6,16'h0066,-16'h0078,-16'h00a3,-16'h0080,16'h00f8,16'h0135,16'h002c,16'h008f,-16'h004a,-16'h0078,16'h01af,-16'h01a6,-16'h014d,16'h0077,16'h0170,16'h002e,-16'h0017,16'h0011,-16'h01ce,16'h00d3,16'h009b,16'h0166,-16'h006c,16'h0016,16'h00fa,16'h0027,16'h0034,16'h00aa,16'h005e,16'h0078,16'h0102,16'h0123,16'h013f,16'h0027,16'h00a2,16'h0079,-16'h0092,16'h017e,16'h00af,-16'h0050,-16'h00da,-16'h0084,16'h01ee,16'h00da,16'h01a5,16'h00bf,16'h010b,16'h00d0,-16'h00ee,-16'h003e,16'h0096,16'h0002,16'h0103,16'h00b4,16'h004c,16'h0096,16'h009e,16'h000d,16'h003c,16'h0029,16'h0056,16'h0062,16'h00fe,16'h0104,16'h003f,-16'h0073,-16'h0058,-16'h0130,16'h00d1,16'h0103,16'h0072,16'h0055,-16'h0057,-16'h0035,16'h01d8,-16'h00a3,-16'h0033,16'h0174,16'h017d,-16'h0027,-16'h0066,16'h0049,-16'h01f5,16'h006a,16'h00f9,16'h0185,16'h004a,-16'h001c,16'h0177,16'h0004,16'h0009,16'h00b6,16'h007f,16'h00c2,16'h00c3,16'h00fa,16'h00e3,16'h00a7,16'h00a7,16'h0076,-16'h005a,16'h0145,-16'h0033,-16'h0012,-16'h002e,-16'h0038,-16'h00a0,16'h0086,16'h01b4,16'h0082,16'h01a1,16'h014a,-16'h00d5,-16'h0061,16'h0087,16'h002e,16'h0171,16'h00a8,16'h006b,16'h0038,16'h005d,16'h0005,-16'h0017,-16'h0031,-16'h001f,16'h00a0,16'h01c9,16'h00be,-16'h0052,16'h002a,-16'h0026,-16'h0184,16'h00a9,16'h00e7,16'h0057,16'h00ef,-16'h0006,16'h0047,16'h020c,16'h0005,16'h002d,16'h01a1,16'h0176,-16'h010b,-16'h0111,16'h00aa,-16'h018d,16'h009f,16'h010e,16'h00b3,16'h0093,16'h000e,16'h00e6,16'h007b,-16'h001f,16'h00c3,16'h0079,16'h00b2,16'h00a0,16'h00ea,16'h0103,16'h0085,16'h006b,16'h0069,-16'h0076,16'h017e,-16'h0040,16'h0010,-16'h0052,-16'h0025,-16'h01b1,16'h00ec,16'h01b0,16'h002c,16'h0189,16'h016f,-16'h0080,-16'h0007,16'h005d,16'h008c,16'h019d,16'h0056,16'h009e,16'h00b0,-16'h0021,-16'h0040,-16'h0009,-16'h002e,-16'h004c,16'h0027,16'h0120,16'h009a,-16'h0022,-16'h000a,16'h0059,-16'h0122,16'h00f9,16'h00c1,16'h009e,16'h002d,-16'h0072,16'h0050,16'h0161,16'h0102,16'h0029,16'h01f1,16'h0135,-16'h00b6,-16'h00bc,-16'h006a,-16'h019a,16'h0036,16'h0079,-16'h004f,16'h00bd,16'h0028,16'h0087,16'h0047,-16'h0139,16'h0040,16'h0010,16'h00d5,16'h0076,16'h0140,16'h002d,16'h0048,16'h001b,16'h0107,16'h0035,16'h01b5,-16'h001f,16'h0053,16'h003b,-16'h000d,-16'h029a,16'h013a,16'h01ab,16'h007e,16'h01b9,16'h0121,-16'h0041,-16'h0159,16'h00ea,16'h0053,16'h0166,16'h00f3,16'h0070,16'h006e,16'h007a,16'h0046,16'h003d,-16'h00b7,16'h0059,16'h0033,16'h0091,16'h00e0,-16'h004c,16'h009e,-16'h001f,-16'h0026,16'h0174,16'h0122,16'h004c,16'h008e,-16'h0072,16'h0084,16'h003e,16'h011f,-16'h006b,16'h0208,16'h01d3,16'h0050,16'h004e,-16'h00e6,-16'h0132,-16'h005e,-16'h0036,-16'h0026,16'h0074,16'h0035,-16'h002d,16'h0040,-16'h010a,16'h00c3,16'h006a,16'h0103,16'h0091,16'h0087,-16'h0009,-16'h0075,-16'h0011,16'h00f7,16'h00ae,16'h019f,-16'h0037,16'h005b,-16'h001a,16'h0007,-16'h016e,16'h00dd,16'h0189,16'h008f,16'h0198,16'h0125,-16'h0037,-16'h01c0,16'h012f,-16'h0006,16'h016e,16'h006e,16'h007f,16'h0047,16'h00be,-16'h000d,16'h004c,-16'h00af,16'h00fa,16'h0084,16'h002f,16'h010b,-16'h0045,16'h0049,-16'h0001,-16'h0092,16'h01ae,16'h00c4,-16'h002f,16'h003b,-16'h0081,16'h00d8,-16'h0010,16'h012d,-16'h003d,16'h019e,16'h01b8,16'h0017,16'h00ad,-16'h0146,-16'h009b,16'h0009,-16'h005a,-16'h0106,-16'h0012,16'h0090,16'h0016,-16'h0033,-16'h00e4,16'h0097,16'h010a,16'h00c1,16'h015a,16'h0045,16'h007a,-16'h0072,-16'h001a,16'h00b3,16'h0093,16'h01fe,-16'h00b4,-16'h0014,16'h0029,16'h0060,-16'h0006,16'h00d4,16'h01bc,-16'h0016,16'h01e6,16'h00c7,-16'h0033,-16'h014b,16'h0114,16'h002f,16'h0177,16'h0024,16'h00c7,16'h0070,16'h00db,-16'h009b,16'h0114,-16'h00c4,16'h004b,16'h006c,16'h000c,16'h00ab,-16'h0034,16'h00c9,16'h00c5,-16'h0065,16'h0180,16'h008b,-16'h000d,16'h00c5,16'h0096,16'h00ac,16'h0019,16'h012b,-16'h0079,16'h00f0,16'h01d0,-16'h0076,16'h010d,-16'h00f1,16'h0004,16'h008a,16'h0017,-16'h007d,-16'h0085,16'h0025,-16'h000b,16'h0002,-16'h0076,16'h00a8,16'h0132,16'h00c6,16'h0131,16'h009f,16'h00dd,16'h0009,16'h00d1,16'h0068,-16'h0008,16'h01f0,-16'h00a2,-16'h000c,16'h007b,-16'h007f,16'h008b,16'h0111,16'h01a7,-16'h006f,16'h01b1,16'h0067,-16'h0035,-16'h00c0,16'h00c7,-16'h0005,16'h00bf,-16'h0004,16'h0078,16'h008b,16'h0099,-16'h00e9,16'h00dd,-16'h020f,16'h0025,16'h004b,-16'h0011,16'h00d1,-16'h006b,16'h00b0,16'h00ee,-16'h0032,16'h0169,16'h008e,-16'h0005,16'h017e,16'h009d,16'h00dc,-16'h00b4,16'h0111,-16'h0091,-16'h032d,16'h01a8,-16'h007d,16'h01f8,-16'h006e,16'h00a9,16'h00b3,16'h000f,16'h00a7,-16'h00c4,16'h003f,-16'h001f,-16'h0094,-16'h0060,16'h0065,16'h0127,16'h006b,16'h00ed,16'h0158,16'h0080,16'h0018,16'h0017,16'h0075,-16'h0002,16'h0164,-16'h0059,-16'h004e,16'h000d,-16'h00b6,16'h00ab,16'h00ad,16'h00b3,-16'h00f5,16'h01f0,16'h001b,-16'h006b,-16'h0001,16'h00f7,-16'h0099,-16'h0099,16'h0034,16'h0056,16'h00c3,16'h004c,-16'h012a,16'h0024,-16'h03fb,-16'h0048,16'h0099,-16'h0100,16'h00f5,-16'h0045,16'h003f,-16'h0031,16'h002e,16'h0143,16'h0083,16'h00bf,16'h0154,16'h00c7,16'h00b7,-16'h0084,16'h00fd,-16'h00f5,-16'h08e7,16'h0176,-16'h008b,16'h01a8,16'h00e6,16'h00da,16'h00f9,-16'h0063,16'h0120,-16'h0100,16'h0047,-16'h0074,-16'h00bb,16'h0058,16'h0147,16'h0127,16'h014a,16'h00cb,16'h00ec,-16'h007c,16'h008b,-16'h006d,16'h00ea,16'h0052,16'h0170,-16'h0034,-16'h0088,-16'h003e,-16'h0174,16'h0003,16'h00c6,16'h00b8,-16'h00c8,16'h0053,-16'h0087,16'h0040,16'h0067,16'h0105,-16'h00a2,-16'h0080,-16'h002b,16'h00fc,16'h009e,-16'h002c,-16'h00c3,16'h007a,-16'h069d,16'h0069,16'h0072,16'h0016,16'h00d5,16'h0035,-16'h0052,16'h006f,-16'h0017,16'h00e4,-16'h0006,16'h0066,-16'h0125,16'h00a2,-16'h00a3,-16'h00a2,16'h0075,-16'h01e5,-16'h0a2f,16'h0123,-16'h0016,16'h01c9,16'h003f,16'h00c4,16'h007f,-16'h0028,16'h016e,-16'h00f5,-16'h0037,16'h0045,-16'h0080,16'h009d,16'h0107,16'h014a,16'h00ff,16'h00c2,16'h00c6,-16'h00bf,-16'h000c,-16'h001b,16'h0071,-16'h0057,16'h01c5,-16'h007a,-16'h00e5,-16'h0066,-16'h0185,16'h000b,16'h008e,16'h0047,-16'h002c,-16'h0434,-16'h0070,16'h0007,-16'h0018,16'h00a2,-16'h00b0,16'h0038,-16'h005f,16'h0068,16'h0118,-16'h00ba,-16'h00f7,16'h006b,-16'h06da,16'h005e,16'h00b8,16'h0087,16'h0014,16'h00c8,-16'h003e,16'h001f,-16'h00e9,16'h0149,-16'h001e,-16'h001b,-16'h02e6,16'h00c5,-16'h0231,-16'h0108,-16'h0125,-16'h00dc,-16'h059d,16'h0128,-16'h001d,16'h0172,-16'h00f0,16'h00a6,16'h007b,-16'h00ac,16'h019e,-16'h0097,-16'h00d4,16'h00b5,-16'h0067,16'h0094,16'h00d2,16'h0045,16'h015b,16'h0141,16'h0049,-16'h00f5,16'h00e2,16'h0047,16'h0067,-16'h0011,16'h010c,-16'h0061,16'h002f,-16'h00c3,-16'h006c,16'h00e9,16'h00f2,16'h0049,16'h0018,-16'h088a,16'h0094,-16'h002b,-16'h00a9,16'h0036,-16'h010e,16'h00a7,-16'h009a,16'h0077,16'h00ee,-16'h00e5,-16'h0112,16'h017c,-16'h05bd,16'h0120,16'h01c9,16'h015c,16'h00af,16'h00a8,-16'h0082,-16'h00b6,-16'h010a,16'h00de,16'h0044,16'h000d,-16'h024e,-16'h0037,-16'h0347,-16'h0172,-16'h0134,-16'h008a,-16'h0315,16'h00eb,16'h0008,-16'h0338,-16'h00ec,-16'h0032,16'h001a,-16'h0154,16'h01c5,16'h0059,-16'h002b,16'h0122,-16'h00f2,16'h0095,-16'h0036,16'h0005,16'h0196,16'h0159,16'h00b1,-16'h01d5,16'h00fb,16'h0021,16'h0059,16'h00ac,16'h0077,-16'h0001,16'h003a,-16'h0010,-16'h001e,16'h007a,16'h0043,16'h0041,16'h00e7,-16'h0670,16'h00ec,-16'h008d,-16'h00d3,16'h0047,-16'h00c1,16'h011e,-16'h00dd,16'h0062,-16'h001b,-16'h00ab,-16'h00e6,-16'h0004,-16'h03dc,16'h0158,16'h0294,16'h017e,16'h004a,16'h00c5,-16'h00bb,-16'h0092,-16'h0065,16'h0160,16'h0057,-16'h005d,-16'h01f8,-16'h00ae,-16'h036e,-16'h00d9,-16'h0065,-16'h0113,-16'h018a,16'h0150,-16'h0057,-16'h06f8,-16'h0097,-16'h018f,16'h0093,-16'h00f9,16'h00cc,16'h00dc,16'h0002,16'h00a1,-16'h00c7,16'h0092,16'h002d,-16'h000a,16'h0261,16'h0159,16'h007b,-16'h0273,16'h0050,-16'h0052,-16'h0024,16'h011b,16'h005a,16'h0019,-16'h0013,16'h0096,-16'h000c,16'h002f,-16'h0017,16'h007b,16'h00a7,-16'h032c,16'h007d,16'h0037,-16'h0152,16'h00d8,-16'h006d,16'h011e,-16'h004d,16'h00e1,-16'h0200,16'h0015,-16'h0100,-16'h0151,-16'h034b,16'h00f7,16'h023b,16'h00f3,16'h002f,16'h00c2,16'h0003,-16'h00d2,16'h001e,16'h0148,16'h0024,16'h007f,-16'h00e8,-16'h0151,-16'h02a9,-16'h0153,-16'h0026,-16'h0086,-16'h005e,16'h00f8,-16'h000b,-16'h0617,-16'h0017,-16'h020a,-16'h0024,-16'h0042,16'h00e6,16'h006f,16'h00ac,16'h0015,-16'h0001,16'h0049,16'h0035,-16'h0017,16'h021a,16'h0174,16'h0032,-16'h0263,-16'h0039,-16'h006e,16'h003e,16'h01e1,16'h0024,16'h00d9,16'h0034,16'h0120,16'h0093,16'h002f,16'h0056,16'h0086,16'h0090,-16'h0136,-16'h0098,-16'h0006,-16'h0044,16'h00f0,16'h000f,16'h00f2,-16'h007a,16'h00ac,-16'h0246,-16'h0092,-16'h00f4,-16'h00d8,-16'h02cf,16'h0000,16'h0146,16'h0103,16'h0028,16'h017a,16'h009e,-16'h0114,16'h002c,16'h010e,16'h004a,16'h0068,-16'h006b,-16'h01ce,-16'h01ca,-16'h0120,16'h0020,-16'h0139,16'h00be,16'h01d3,16'h0040,-16'h043c,-16'h0053,-16'h02c3,16'h0128,-16'h0085,16'h006a,16'h0028,16'h0117,16'h004c,16'h008f,16'h0017,16'h0010,16'h009e,16'h0199,16'h0284,-16'h008f,-16'h024d,-16'h0029,-16'h0067,-16'h0053,16'h00d4,16'h00c9,16'h007b,16'h005b,16'h01b7,16'h001d,16'h0003,16'h0089,16'h008c,16'h00e0,-16'h007d,-16'h0244,-16'h009a,16'h0074,16'h0167,16'h0087,16'h016f,16'h011e,-16'h005c,-16'h0051,16'h00f7,16'h0107,16'h0105,16'h013c,-16'h004b,16'h03b1,-16'h0102,16'h01fe,16'h0061,16'h001f,16'h0052,16'h0002,-16'h0078,16'h007d,-16'h00b8,-16'h0121,16'h0022,16'h0258,16'h0025,-16'h004e,-16'h01fc,-16'h00c5,-16'h00ac,-16'h00f3,16'h0070,16'h0377,16'h01ec,16'h00d8,16'h00ac,-16'h0165,-16'h0074,16'h00df,-16'h0055,-16'h0053,16'h026d,-16'h0025,16'h0093,16'h0168,16'h005a,-16'h0018,-16'h0038,16'h006e,-16'h000f,16'h011d,-16'h00ea,16'h00f0,-16'h008b,-16'h0055,16'h0082,-16'h0128,16'h00a5,16'h005c,-16'h011f,-16'h0071,-16'h0087,-16'h000f,-16'h00a3,16'h0140,16'h0083,16'h0041,16'h0159,16'h01e2,-16'h0084,-16'h00cd,16'h0081,16'h012a,16'h0048,16'h013b,16'h00af,16'h0290,-16'h0166,16'h0201,16'h0067,16'h004a,16'h0064,16'h0095,-16'h00a9,16'h004d,-16'h00f6,-16'h0090,16'h0046,16'h000c,16'h00a6,-16'h006b,-16'h02e0,-16'h00b7,-16'h00b8,-16'h00a3,-16'h005f,16'h02ed,16'h0238,16'h0119,16'h0102,-16'h01d3,-16'h00a7,-16'h0039,-16'h007c,16'h00a6,16'h028c,-16'h0008,16'h004c,16'h0089,16'h0123,-16'h000c,-16'h0033,16'h0070,-16'h00b5,16'h00b4,-16'h00d6,16'h0057,-16'h00a0,-16'h0088,16'h00c2,16'h0000,16'h01bc,-16'h0021,-16'h005b,16'h0023,-16'h0071,-16'h0009,-16'h005d,16'h0087,16'h00b5,16'h0092,16'h015a,16'h01c9,-16'h014d,-16'h006e,16'h002f,16'h0039,-16'h0077,16'h0108,16'h0104,16'h01ed,-16'h01a8,16'h0126,16'h004b,16'h0099,-16'h000e,16'h00e0,16'h000f,16'h008f,-16'h009c,-16'h006d,-16'h0073,-16'h000e,16'h01bc,-16'h006c,-16'h0427,-16'h002b,-16'h0070,-16'h013e,-16'h009e,16'h01ce,16'h0112,16'h00a2,16'h005d,-16'h006a,16'h0007,-16'h013d,-16'h0044,16'h0060,16'h01eb,-16'h0003,-16'h0063,16'h00c9,16'h013d,16'h0077,-16'h002e,16'h0080,-16'h00c5,16'h003d,-16'h011c,16'h0078,16'h0048,-16'h00e0,16'h00c6,16'h0070,16'h01f6,-16'h0060,-16'h00cc,-16'h00f1,-16'h0045,16'h0005,-16'h0104,16'h0075,16'h0121,16'h0097,16'h0184,16'h0134,-16'h0212,16'h001e,16'h0043,16'h0017,-16'h005f,16'h0045,16'h00b6,16'h00cb,-16'h0269,16'h00a4,-16'h0118,16'h005a,-16'h003c,16'h000f,-16'h001d,16'h00b6,-16'h00b8,16'h0055,-16'h01ab,-16'h0054,16'h020c,-16'h003d,-16'h03d1,16'h0025,-16'h009e,-16'h00b6,-16'h00ab,16'h01d8,-16'h005d,16'h009d,-16'h0088,16'h00a6,16'h005d,-16'h0109,-16'h00ba,16'h00ac,16'h010c,16'h003d,-16'h005a,16'h011b,16'h01a2,16'h0042,-16'h000c,16'h0086,16'h002d,16'h0078,-16'h006c,16'h00d5,16'h0028,-16'h00c8,16'h0185,16'h0224,16'h0181,-16'h00a5,-16'h00d9,-16'h00b9,16'h0069,-16'h0006,-16'h0143,16'h0068,16'h00cd,16'h008c,16'h01b7,16'h00af,-16'h01bb,16'h002f,-16'h002a,16'h0069,16'h0008,-16'h001a,16'h00bb,16'h00ab,-16'h02c2,16'h0019,-16'h00a5,16'h000b,16'h002d,-16'h0016,16'h005b,16'h012f,-16'h00db,16'h0096,-16'h0274,-16'h0037,16'h01e1,16'h0051,-16'h023a,16'h0075,-16'h009e,-16'h0001,-16'h0058,16'h0187,16'h000c,16'h004f,-16'h0225,16'h01c2,16'h0075,-16'h0159,-16'h008f,16'h0100,16'h013e,-16'h0049,16'h0030,16'h0064,16'h0222,16'h0040,16'h0071,16'h00ab,16'h00d7,16'h00a4,-16'h0010,16'h0163,16'h0069,-16'h0046,16'h008e,16'h0215,16'h0062,-16'h00c3,-16'h0137,-16'h00cf,16'h0056,16'h0080,-16'h01df,16'h0060,16'h00c8,16'h0028,16'h0128,16'h0174,-16'h01e1,16'h00d7,16'h001a,16'h0024,16'h0073,-16'h0010,16'h00e4,16'h00f7,-16'h0288,16'h00a0,-16'h002a,-16'h008c,-16'h003a,-16'h0076,16'h000a,16'h010f,-16'h00c4,16'h00d8,-16'h021d,16'h0090,16'h0226,16'h0172,-16'h015c,16'h0100,-16'h0047,-16'h0054,-16'h000f,16'h01d6,-16'h0004,16'h0092,-16'h01f4,16'h01c1,-16'h009e,-16'h019a,-16'h00f7,16'h004d,16'h00ee,-16'h00da,16'h0068,-16'h0044,16'h0206,16'h006f,-16'h0003,16'h00e4,16'h009d,16'h0035,-16'h0097,16'h0180,16'h00d6,16'h001a,16'h00a0,16'h0205,-16'h005a,-16'h0066,-16'h0111,-16'h00fd,16'h0128,16'h0030,-16'h01ed,16'h0065,16'h0131,16'h005a,16'h014a,16'h00dd,-16'h016a,16'h0098,16'h006a,16'h0097,16'h017a,-16'h0057,16'h0051,16'h0110,-16'h025a,16'h012b,16'h0047,-16'h004f,-16'h000f,-16'h0092,16'h0083,16'h01a6,-16'h0056,16'h00ca,-16'h00c2,16'h008a,16'h02c1,16'h01e3,-16'h01ec,16'h00f1,-16'h0040,-16'h0088,16'h0081,16'h0179,16'h0059,16'h00db,-16'h00a9,16'h011f,-16'h018e,-16'h00c4,16'h0016,16'h0034,-16'h00bb,-16'h000e,-16'h002e,-16'h0085,16'h0187,16'h0026,-16'h0094,16'h00ac,16'h0042,16'h006c,-16'h00d6,16'h0169,16'h0088,16'h0056,16'h00a6,16'h0249,-16'h012d,-16'h0030,-16'h017b,-16'h00c4,16'h0035,16'h00c1,-16'h0194,16'h00ad,16'h005a,16'h0055,16'h0146,16'h0142,-16'h028e,16'h0034,16'h0036,16'h001d,16'h015a,-16'h0015,16'h007a,16'h0109,-16'h00ee,16'h00fd,-16'h001e,16'h006f,16'h004e,-16'h00c6,16'h00c0,16'h00f9,-16'h00aa,16'h0033,16'h0031,16'h00b1,16'h0241,16'h0189,-16'h01b6,16'h009a,-16'h001a,-16'h023e,16'h008a,16'h0263,16'h01e7,16'h0141,16'h006f,-16'h000d,-16'h0157,-16'h00ef,16'h00cd,-16'h000b,-16'h014f,16'h0044,-16'h017f,-16'h0011,16'h00e4,-16'h0006,-16'h0065,16'h00cb,16'h0067,16'h00d7,-16'h016e,16'h018c,16'h0002,16'h009f,16'h0059,16'h0235,-16'h01f2,16'h0037,-16'h01b3,-16'h001d,16'h00ae,16'h013f,-16'h01b2,-16'h0009,16'h00a1,16'h0016,16'h00fa,16'h0153,-16'h024c,-16'h0022,16'h0152,16'h009a,16'h00a9,16'h0045,16'h0092,16'h0127,16'h0043,16'h0163,-16'h0026,16'h0108,-16'h0028,-16'h00b5,16'h00bb,16'h00ed,16'h004b,-16'h00ca,16'h0115,16'h00e1,16'h021b,16'h00f8,-16'h014f,16'h0059,-16'h001c,-16'h028f,-16'h0026,16'h0134,16'h01c3,16'h00f9,16'h0037,-16'h010f,-16'h0055,-16'h00a6,16'h0146,16'h002f,-16'h00af,16'h01b4,-16'h019d,-16'h0086,16'h0194,16'h00e8,16'h0010,16'h0096,16'h00ed,16'h0056,-16'h013c,16'h0139,-16'h0018,16'h00c3,-16'h0060,16'h01fb,-16'h01f2,16'h0080,-16'h019c,16'h0029,16'h0043,16'h017d,-16'h0206,-16'h002a,16'h0095,-16'h0019,16'h0134,16'h0094,-16'h01b9,-16'h0007,16'h014c,16'h00f0,16'h005c,16'h0078,-16'h002d,16'h013b,16'h00ba,16'h01b0,-16'h00db,16'h00dd,-16'h001b,-16'h0116,16'h00de,16'h00bc,16'h0076,-16'h008c,16'h0142,16'h0154,16'h020c,-16'h00e8,-16'h012d,16'h0075,16'h0059,-16'h0129,16'h00a1,-16'h00cc,16'h0167,16'h00bc,16'h0067,-16'h0072,16'h0135,-16'h0038,-16'h0158,16'h0006,-16'h0021,16'h014b,-16'h016c,-16'h00cf,16'h01b9,16'h00be,16'h010b,16'h0097,16'h00b2,16'h0068,-16'h00ec,16'h0163,-16'h004a,16'h0112,-16'h016f,16'h012f,-16'h00f7,16'h007b,-16'h009d,16'h0038,16'h00b9,16'h01e0,-16'h01b4,-16'h00ac,16'h00c1,-16'h0038,16'h0174,16'h00ec,-16'h010d,16'h00b9,16'h00d3,16'h0097,-16'h000f,16'h005e,16'h003c,16'h00fc,16'h0122,16'h010f,-16'h00ac,16'h013c,-16'h0089,-16'h00c5,16'h0121,16'h0032,16'h008e,-16'h0082,16'h01a6,16'h007e,16'h0120,-16'h0235,-16'h018d,16'h002c,16'h0080,16'h00b7,16'h00b6,-16'h0230,16'h009b,16'h010c,16'h00bc,-16'h0076,16'h00ea,-16'h0011,-16'h02fc,-16'h0014,-16'h007d,16'h00f3,-16'h005c,-16'h00df,16'h015d,16'h0113,16'h012f,16'h007e,16'h00b4,-16'h0042,-16'h007a,16'h01bf,16'h0092,16'h00c5,-16'h00b4,16'h00a5,16'h0094,16'h004d,16'h0055,16'h0042,16'h00c2,16'h0156,-16'h015e,-16'h00a0,16'h0110,-16'h002d,16'h00f9,16'h0133,-16'h00a1,16'h008f,16'h011f,16'h00d5,16'h0027,16'h0093,16'h0028,16'h007c,16'h0155,16'h011a,-16'h0097,16'h005d,-16'h007d,-16'h00a1,16'h0138,16'h004f,16'h0025,-16'h001b,16'h0107,-16'h00a2,16'h0172,-16'h0279,-16'h0196,16'h0014,16'h0054,16'h01d6,16'h00a1,-16'h02a6,-16'h0070,16'h0140,16'h0027,16'h010e,16'h0050,-16'h0023,-16'h02d8,16'h0013,-16'h0021,16'h0054,-16'h000b,-16'h002a,16'h0147,16'h00da,16'h00e2,16'h00a3,16'h0113,16'h0012,-16'h00ad,16'h022f,16'h0062,-16'h0044,-16'h0165,16'h0032,16'h01b0,16'h002f,16'h0034,16'h00fa,16'h002c,16'h0108,-16'h0177,-16'h0193,16'h00cb,-16'h0002,16'h00c2,16'h00ca,-16'h012d,16'h004e,16'h007e,16'h0041,16'h00d5,16'h0034,16'h0050,16'h005a,16'h00e1,16'h0142,-16'h004d,-16'h0026,-16'h00b1,-16'h0007,16'h010f,16'h0072,16'h0008,16'h011d,-16'h0008,-16'h008f,16'h01db,-16'h01a6,-16'h0171,-16'h002c,16'h00d1,16'h00eb,-16'h0009,-16'h023e,-16'h01ea,16'h00dc,16'h0041,16'h017f,16'h0031,16'h000b,-16'h0152,-16'h0098,16'h0020,16'h008c,16'h0076,16'h003b,16'h0090,16'h00b9,16'h00f9,16'h00b8,16'h009a,-16'h0052,-16'h00f8,16'h01f9,16'h00e7,-16'h000e,-16'h0164,-16'h000e,16'h0260,16'h001a,16'h001d,16'h00e6,16'h0036,16'h007b,-16'h0179,-16'h0163,16'h0135,16'h0008,16'h00a9,16'h00fb,-16'h0114,16'h006f,16'h00d0,-16'h0046,16'h00a7,16'h0034,16'h0076,16'h006f,16'h00d0,16'h0147,16'h0026,-16'h0059,-16'h0069,-16'h003f,16'h0114,16'h00cb,16'h0029,16'h0120,-16'h0094,-16'h00ad,16'h0178,-16'h0122,-16'h0189,16'h006a,16'h00ee,16'h00da,-16'h0027,-16'h016c,-16'h01d4,16'h00f7,16'h00db,16'h012a,16'h006c,16'h0063,16'h00f3,-16'h00ce,16'h005c,16'h007e,16'h000a,16'h00ad,16'h006d,16'h0180,16'h0158,16'h00e4,16'h00b7,-16'h0020,-16'h00f7,16'h01d3,16'h00ad,16'h004a,-16'h0157,-16'h0006,16'h0180,16'h000f,16'h010f,16'h00ca,16'h0054,16'h00ad,-16'h01f7,-16'h0120,16'h006b,16'h0023,16'h010b,16'h0103,-16'h00d4,16'h003b,16'h006f,-16'h0052,16'h0040,16'h0000,16'h005a,16'h00ba,16'h0129,16'h012e,-16'h000a,-16'h0098,-16'h000a,-16'h0084,16'h00b6,16'h00f2,16'h00df,16'h00f4,-16'h0077,-16'h0011,16'h01aa,16'h005e,-16'h00fa,16'h0140,16'h0179,16'h0036,16'h0016,-16'h003d,-16'h01b0,16'h00e8,16'h0157,16'h0003,16'h0102,-16'h0034,16'h017a,-16'h0099,16'h0016,16'h008a,16'h0014,16'h00ab,16'h002f,16'h0114,16'h00ea,16'h011c,16'h0049,16'h0054,-16'h0063,16'h01cf,16'h006b,-16'h0053,-16'h009b,-16'h00cd,-16'h0095,-16'h0045,16'h01b5,16'h00df,16'h00a3,16'h00ca,-16'h017e,-16'h012c,16'h007e,16'h0010,16'h0163,16'h00bf,-16'h00e7,16'h00ca,16'h002b,-16'h00d6,-16'h0006,-16'h0038,16'h0008,16'h00cb,16'h0105,16'h01b8,-16'h0072,-16'h0049,-16'h0038,-16'h00e9,16'h00ad,16'h00e1,16'h009d,16'h0106,-16'h0013,-16'h0030,16'h01d5,16'h00eb,16'h002d,16'h018e,16'h01e2,-16'h00ed,-16'h0056,-16'h0014,-16'h0112,16'h00cf,16'h0170,-16'h0005,16'h0053,-16'h004e,16'h00ae,-16'h0006,16'h0035,16'h00b0,16'h0002,16'h010f,16'h001e,16'h012a,16'h00d2,16'h0050,16'h009a,16'h0103,-16'h0089,16'h01bd,16'h0054,16'h010c,-16'h002f,-16'h00c9,-16'h01fa,16'h0001,16'h011b,16'h0098,16'h0059,16'h00ed,-16'h014a,-16'h00c9,16'h00ba,16'h00d0,16'h0208,16'h0111,-16'h017f,16'h0080,16'h0067,-16'h00ba,-16'h0082,-16'h0166,16'h0009,16'h00ad,16'h00a2,16'h0168,-16'h0026,16'h0015,16'h0005,-16'h0061,16'h0126,16'h0079,16'h006e,16'h00c8,-16'h00ab,16'h0025,16'h00e2,16'h0095,16'h0002,16'h024b,16'h017f,-16'h00df,-16'h003d,-16'h00b0,-16'h009f,16'h003f,16'h009f,-16'h00ae,16'h00b0,-16'h005b,16'h007d,-16'h0020,16'h0006,16'h00fb,-16'h0043,16'h00ca,-16'h001d,16'h0057,16'h0002,16'h0048,16'h0062,16'h00f8,-16'h0021,16'h0224,-16'h0033,16'h0128,16'h0076,-16'h00b9,-16'h02c9,16'h00c1,16'h0092,16'h002d,16'h0131,16'h0120,-16'h015d,-16'h00c1,16'h0148,16'h009f,16'h0211,16'h00db,-16'h00a2,16'h004f,16'h0010,-16'h00f7,16'h002d,-16'h0148,-16'h0010,16'h0076,16'h003e,16'h011a,-16'h008c,16'h003d,-16'h004d,-16'h0016,16'h0156,16'h0060,16'h0070,16'h00ba,-16'h00cc,16'h008e,16'h0057,16'h0168,-16'h0099,16'h024b,16'h01c1,16'h0002,16'h007b,-16'h013b,-16'h0030,16'h00bc,16'h0067,-16'h00cf,-16'h0020,-16'h0042,-16'h0004,-16'h0037,16'h0039,16'h00c6,16'h0066,16'h0092,16'h0021,16'h0084,16'h0037,16'h000c,-16'h0035,16'h00c2,-16'h002a,16'h01e3,-16'h004c,16'h00fc,16'h0004,-16'h00b6,-16'h018a,16'h0043,16'h00eb,16'h0059,16'h0113,16'h0137,-16'h019d,-16'h0140,16'h0139,16'h0016,16'h0190,16'h00f9,-16'h00b5,16'h006f,16'h00df,-16'h018d,16'h008e,-16'h01fb,16'h0000,16'h006f,16'h006d,16'h018b,-16'h0034,-16'h0011,-16'h001b,16'h0020,16'h0161,16'h0099,16'h0009,16'h008c,-16'h0011,16'h0155,16'h00da,16'h00e3,-16'h0025,16'h0206,16'h01f8,16'h0006,16'h0138,-16'h00c6,-16'h0007,16'h0085,16'h003b,-16'h003a,-16'h00da,16'h0001,-16'h00a0,16'h001f,-16'h0065,16'h0068,16'h016d,16'h0100,16'h004e,-16'h0027,-16'h0013,16'h00bf,16'h003a,16'h0123,16'h0098,16'h0156,-16'h0044,16'h008a,16'h0049,-16'h00df,16'h0014,16'h001a,16'h0106,-16'h0065,16'h0153,16'h0142,-16'h023d,-16'h00c0,16'h0150,16'h0048,16'h01c7,16'h006d,-16'h0051,16'h000a,16'h00c7,-16'h015f,16'h00f7,-16'h037d,-16'h002d,16'h00bc,16'h0029,16'h017a,-16'h0040,16'h0073,-16'h001c,16'h0009,16'h013b,16'h0026,16'h0005,16'h0065,16'h00a6,16'h00ae,16'h00cd,16'h00cc,-16'h008c,16'h0108,16'h01a5,-16'h002d,16'h0157,-16'h00c1,16'h0075,16'h00b8,-16'h0060,-16'h0002,-16'h00dd,16'h0041,-16'h0036,-16'h005e,-16'h00ef,16'h010c,16'h00e2,16'h00dc,16'h00e0,16'h003f,16'h0036,16'h00c8,-16'h0002,16'h0125,16'h002d,16'h0118,-16'h004a,16'h0016,16'h0098,-16'h00c2,16'h00b0,16'h007f,16'h00fc,-16'h0068,16'h0144,16'h008f,-16'h0285,16'h0028,16'h005a,16'h008a,16'h00f4,16'h0052,16'h0012,16'h0122,16'h0016,-16'h0144,16'h005a,-16'h0591,-16'h0030,16'h00c5,-16'h002d,16'h00e9,16'h0028,16'h00f7,16'h006b,16'h0060,16'h010b,16'h00bd,-16'h0018,16'h018a,16'h0089,16'h004a,16'h0067,16'h00b1,-16'h0015,-16'h02a3,16'h01d1,-16'h0016,16'h0199,-16'h0074,16'h00bc,16'h0153,-16'h0052,16'h0083,-16'h00c0,16'h003c,-16'h0043,-16'h0084,-16'h0002,16'h0078,16'h0067,16'h00f1,16'h0113,16'h00c4,-16'h00ff,16'h00f4,-16'h0038,16'h00a6,-16'h0021,16'h00e3,16'h002b,16'h0006,16'h0006,-16'h00cc,16'h00da,16'h0095,16'h0077,-16'h00cd,16'h0105,16'h006a,-16'h01bf,16'h009e,-16'h002c,16'h0004,16'h0003,-16'h002e,16'h0093,16'h016e,-16'h0047,-16'h00dd,16'h005f,-16'h06f1,-16'h0036,16'h00c7,-16'h0023,16'h00d7,16'h001e,16'h00a5,16'h00bf,16'h0056,16'h00a2,16'h00d0,16'h001f,16'h00cd,16'h00de,-16'h0077,16'h0032,16'h0075,-16'h00e2,-16'h093e,16'h0100,16'h0005,16'h019a,16'h0003,16'h0088,16'h0170,-16'h007a,16'h019e,-16'h00c9,16'h0025,-16'h0078,-16'h0112,16'h0023,16'h004d,16'h0044,16'h00f9,16'h00b9,16'h0107,-16'h0173,16'h00a4,-16'h00c9,16'h00c9,-16'h0099,16'h0201,16'h0052,-16'h006d,-16'h0032,-16'h00e8,16'h0026,16'h0083,16'h00cd,-16'h00fe,-16'h0056,-16'h001a,-16'h0143,16'h0022,16'h007e,-16'h003b,-16'h001c,-16'h0064,16'h003c,16'h015b,-16'h0068,-16'h009b,16'h00ab,-16'h06a0,16'h0087,16'h00c1,-16'h0016,16'h007f,16'h0078,16'h000e,16'h0034,-16'h0092,16'h00c5,16'h0058,16'h00ac,-16'h01d6,16'h0042,-16'h01b1,16'h0039,-16'h00c2,-16'h01b5,-16'h0aa1,16'h0151,-16'h0032,16'h01ec,-16'h003a,16'h005f,16'h00fd,16'h0056,16'h0177,-16'h007f,-16'h000b,16'h004b,-16'h0135,16'h0003,16'h007f,16'h0052,16'h0172,16'h00bd,16'h0092,-16'h0255,16'h0090,-16'h0023,16'h00e0,-16'h003b,16'h01a3,-16'h0028,-16'h0020,-16'h0091,-16'h00d1,-16'h003e,16'h006a,16'h00aa,-16'h007d,-16'h063f,-16'h0039,-16'h016f,-16'h0090,16'h0098,-16'h00f5,16'h00a5,16'h0050,16'h0076,16'h0168,-16'h00e1,-16'h00db,16'h00f2,-16'h0551,16'h00c3,16'h00e0,16'h0000,16'h0012,16'h00b0,-16'h00b2,-16'h000b,-16'h0110,16'h00c5,16'h004c,16'h0023,-16'h0326,16'h001a,-16'h031f,16'h0015,-16'h0191,-16'h00a5,-16'h05a6,16'h0182,16'h0004,16'h014c,-16'h016b,-16'h0050,16'h0094,16'h002b,16'h01b7,-16'h0001,-16'h0091,16'h0134,-16'h0072,16'h006d,16'h0026,16'h002a,16'h0107,16'h0024,16'h004d,-16'h0230,16'h00b0,16'h002a,16'h0040,16'h0035,16'h016c,-16'h0043,16'h006e,-16'h0057,-16'h0035,16'h0019,16'h0057,16'h0118,-16'h002d,-16'h099e,-16'h0004,-16'h00df,-16'h006c,16'h0003,-16'h013d,16'h0106,16'h0043,16'h0076,16'h00fb,-16'h00d1,-16'h00a0,16'h00db,-16'h03ad,16'h0070,16'h01c0,16'h00fb,16'h0017,16'h00e0,-16'h00fe,-16'h00ca,-16'h00a4,16'h009a,16'h007d,-16'h005f,-16'h021f,-16'h002b,-16'h03fa,-16'h003f,-16'h01d6,-16'h0099,-16'h02cd,16'h011e,-16'h001e,-16'h0330,-16'h0188,-16'h0149,16'h00ca,-16'h0073,16'h01bb,-16'h0007,-16'h009c,16'h0127,-16'h0122,16'h008a,16'h0018,-16'h007a,16'h01ba,16'h010f,-16'h0014,-16'h0359,16'h00ad,-16'h005f,16'h0060,16'h00d7,16'h00d8,16'h0038,16'h0028,16'h007c,-16'h003c,16'h00ea,16'h0021,16'h0054,16'h00b9,-16'h0612,16'h0110,-16'h0167,-16'h0099,16'h00f5,-16'h00a8,16'h0196,-16'h0016,16'h0085,16'h0091,-16'h006b,-16'h00bb,-16'h0015,-16'h02f5,16'h00a6,16'h0286,16'h0106,-16'h0055,16'h00e2,-16'h0035,-16'h00ce,16'h0033,16'h013e,-16'h0017,-16'h0005,-16'h01df,-16'h009c,-16'h0303,-16'h001c,-16'h0074,-16'h0096,-16'h016b,16'h01e5,16'h0065,-16'h06b7,-16'h00b5,-16'h025b,16'h0068,-16'h005a,16'h015d,16'h0040,-16'h0012,16'h00a4,-16'h00db,16'h000c,16'h0045,-16'h0056,16'h022f,16'h005f,16'h004c,-16'h038c,16'h001c,-16'h004a,-16'h0015,16'h01b4,16'h0063,16'h00fe,16'h00b2,16'h0111,-16'h0013,16'h00ac,-16'h003b,16'h005c,16'h004e,-16'h02f7,16'h00ca,-16'h012e,-16'h0075,16'h0108,-16'h0094,16'h01a3,16'h005c,16'h004e,-16'h0146,-16'h00b3,-16'h00af,-16'h014d,-16'h0324,16'h001c,16'h0287,16'h0088,-16'h009f,16'h016a,16'h0042,-16'h014e,16'h0054,16'h00af,-16'h001a,16'h0009,-16'h00f4,-16'h00a4,-16'h0250,-16'h0047,-16'h009e,-16'h0063,-16'h004d,16'h018a,-16'h0029,-16'h05e5,-16'h002c,-16'h0222,16'h0001,-16'h007b,16'h0141,16'h0098,16'h008d,16'h0029,-16'h0045,16'h0045,16'h000c,-16'h005c,16'h01b7,16'h010c,-16'h000b,-16'h0211,-16'h00ad,-16'h009b,-16'h003f,16'h0204,16'h00f1,16'h015b,16'h00c7,16'h01a8,16'h007f,16'h008c,-16'h0060,16'h007a,16'h00b1,-16'h00f2,-16'h007a,-16'h0114,16'h004d,16'h001e,-16'h00a4,16'h0129,16'h00a0,16'h0040,-16'h029c,-16'h00f6,-16'h0161,-16'h0186,-16'h025d,16'h001c,16'h0232,16'h010d,16'h004a,16'h00de,16'h00c0,-16'h01a7,16'h009c,16'h0186,16'h0052,16'h0076,-16'h0112,-16'h00f2,-16'h01bc,-16'h0032,-16'h009e,-16'h00ff,16'h00de,16'h01d5,16'h00c8,-16'h044e,-16'h0031,-16'h025a,16'h00bc,-16'h00c9,-16'h0001,16'h0076,16'h018b,16'h001f,16'h00be,16'h00c2,-16'h004c,16'h0132,16'h0131,16'h019a,-16'h0047,-16'h0229,-16'h0021,-16'h0062,-16'h0066,16'h016b,16'h0117,16'h0056,16'h003a,16'h01ae,16'h0048,-16'h001e,-16'h005b,16'h000a,16'h0049,16'h0003,-16'h0105,-16'h00e2,16'h0084,16'h0181,16'h010b,16'h012d,16'h007f,-16'h012e,16'h001e,16'h00f7,16'h0084,16'h0136,16'h01c6,-16'h00e6,16'h02a8,-16'h00e3,16'h0257,16'h0053,-16'h0012,16'h002e,16'h0037,-16'h0041,16'h00ab,-16'h0162,-16'h0063,16'h005d,16'h028b,-16'h001c,-16'h007e,-16'h0253,-16'h0051,-16'h0011,-16'h000b,-16'h0032,16'h03ad,16'h01c1,16'h0138,16'h00d9,-16'h0197,-16'h00ba,16'h00fd,-16'h005f,-16'h0009,16'h0286,-16'h0039,16'h001c,16'h010d,16'h0028,-16'h001c,-16'h000c,16'h0035,16'h009e,16'h00dc,-16'h0091,16'h0165,-16'h0098,-16'h0035,16'h009f,-16'h00ff,16'h00f2,16'h0033,-16'h0104,-16'h010d,-16'h00e8,16'h010d,-16'h0067,16'h015b,16'h0171,16'h0096,16'h00b4,16'h01ae,-16'h0115,-16'h0086,16'h00aa,16'h0047,16'h00c7,16'h0129,16'h0087,16'h02c8,-16'h0200,16'h01b1,16'h0032,-16'h0033,16'h0019,16'h00d5,-16'h0088,16'h0104,-16'h00ec,-16'h00bc,16'h0064,16'h00a1,16'h004e,-16'h0028,-16'h030d,16'h0007,-16'h0058,-16'h0082,16'h0021,16'h0354,16'h01d5,16'h012e,16'h0057,-16'h0155,-16'h00fe,16'h0053,-16'h0098,16'h0034,16'h0236,16'h0001,16'h000e,16'h0169,16'h00e5,-16'h0026,16'h005a,16'h001c,-16'h0061,16'h00c9,-16'h0072,16'h00c5,16'h0041,16'h002d,16'h0158,-16'h0001,16'h0154,-16'h006a,-16'h017e,-16'h00a0,-16'h004c,16'h0089,-16'h0092,16'h0089,16'h00f2,16'h009e,16'h015b,16'h01cf,-16'h0189,16'h0057,16'h0052,-16'h0024,16'h003d,16'h00a7,16'h013b,16'h023a,-16'h0161,16'h00c0,16'h0000,16'h0092,-16'h0001,16'h00b2,-16'h00f0,16'h009d,-16'h00be,-16'h002c,-16'h007b,-16'h000c,16'h0074,16'h0027,-16'h03b0,-16'h0044,-16'h0065,-16'h00a3,-16'h0079,16'h0350,16'h017b,16'h00ed,16'h000f,-16'h0144,-16'h0038,-16'h008a,-16'h0127,16'h0032,16'h022e,-16'h00a4,-16'h0065,16'h017d,16'h00e9,-16'h004f,16'h0015,16'h00bf,-16'h003f,16'h0034,-16'h011c,16'h00ab,-16'h002c,-16'h006c,16'h014e,16'h00c6,16'h01e0,-16'h0017,-16'h011e,-16'h00c6,16'h001f,16'h0052,-16'h00b4,16'h00e0,16'h00b3,16'h00a0,16'h01c2,16'h01da,-16'h027c,16'h0065,16'h0058,-16'h0070,-16'h0004,16'h0051,16'h0142,16'h018c,-16'h0256,16'h0048,-16'h008d,16'h00c6,-16'h0078,16'h00b9,-16'h0128,16'h003f,-16'h0057,-16'h0052,-16'h01e9,-16'h0047,16'h0164,16'h00ab,-16'h0358,-16'h000c,-16'h0103,-16'h0026,-16'h0084,16'h0224,16'h00d0,16'h0068,-16'h00b0,-16'h0035,16'h0093,-16'h01b3,-16'h00ce,-16'h004f,16'h017a,-16'h00f2,16'h0045,16'h0127,16'h012a,-16'h0069,-16'h004a,16'h0086,16'h0067,16'h003e,-16'h00b0,16'h00a2,16'h0079,-16'h00cd,16'h0117,16'h021b,16'h0183,-16'h0030,-16'h00fb,-16'h00e2,16'h004e,16'h0069,-16'h00b7,16'h00f9,16'h00ec,16'h00ae,16'h0129,16'h018f,-16'h036f,16'h013c,16'h00aa,16'h003d,16'h0072,16'h0047,16'h0168,16'h00ce,-16'h0264,-16'h0021,-16'h00db,-16'h0046,-16'h008d,16'h001c,-16'h0098,16'h0043,-16'h0078,16'h0078,-16'h02b6,16'h0018,16'h01ed,16'h00e7,-16'h01a3,16'h0114,-16'h00f4,16'h0001,-16'h0057,16'h01cd,16'h006d,16'h00b5,-16'h01ab,16'h0156,16'h003d,-16'h01dd,-16'h00de,-16'h000d,16'h01dc,-16'h0079,16'h0035,16'h008b,16'h0182,16'h007b,-16'h0048,16'h00e9,16'h006d,16'h00a1,-16'h010c,16'h00b3,-16'h0020,-16'h0085,16'h0133,16'h01dc,16'h00ad,-16'h012e,-16'h0130,-16'h0103,16'h0060,16'h0033,-16'h01aa,16'h00b8,16'h006c,16'h0065,16'h0177,16'h01c6,-16'h02d6,16'h01a6,16'h0095,16'h005b,16'h005e,-16'h001a,16'h0172,16'h0051,-16'h019f,16'h000a,16'h00a2,-16'h0113,-16'h002d,-16'h0034,-16'h0064,16'h005e,-16'h00bf,16'h0127,-16'h01f7,16'h0069,16'h0271,16'h0158,-16'h00fe,16'h0081,-16'h0116,16'h000b,-16'h0040,16'h022c,16'h0051,16'h009d,-16'h0142,16'h01af,-16'h0082,-16'h0210,-16'h00d9,-16'h0042,16'h00e5,-16'h013a,16'h000f,16'h0060,16'h018f,-16'h0008,-16'h00a0,16'h00cf,16'h0052,16'h0047,-16'h008f,16'h0067,-16'h0019,16'h001f,16'h00e3,16'h01fb,-16'h0013,-16'h019d,-16'h0194,-16'h011a,16'h0041,16'h00b1,-16'h013d,16'h010d,16'h0084,-16'h002e,16'h0108,16'h01b7,-16'h02cf,16'h012a,16'h00c7,16'h00a8,16'h00ec,16'h0000,16'h016b,16'h0065,-16'h013a,16'h0092,16'h0088,16'h0004,16'h0046,16'h0011,-16'h0011,-16'h0049,-16'h009a,16'h00d7,-16'h008e,16'h0104,16'h02e6,16'h01df,-16'h013d,16'h010a,-16'h012e,-16'h0090,16'h0065,16'h0221,16'h00b8,16'h010b,-16'h00ca,16'h00f7,-16'h018b,-16'h0181,-16'h0015,-16'h0079,16'h001c,-16'h00ba,-16'h00d1,-16'h0019,16'h01dc,-16'h0008,-16'h0081,16'h0124,16'h00a5,16'h0080,-16'h008d,16'h0128,-16'h0025,-16'h0016,16'h00a4,16'h0158,-16'h0131,-16'h011b,-16'h01dc,-16'h010d,-16'h0034,16'h007b,-16'h0182,16'h0091,16'h00b1,16'h002e,16'h0146,16'h0146,-16'h0343,16'h00fb,16'h012c,16'h00d4,16'h0093,16'h0062,16'h0180,16'h00b5,-16'h0067,16'h00d5,16'h0046,16'h0016,16'h0024,16'h0024,16'h0064,-16'h0061,-16'h0026,16'h00ab,-16'h0003,16'h00f8,16'h0278,16'h01a4,-16'h0170,16'h0116,-16'h00a6,-16'h01a6,16'h0084,16'h01ea,16'h017a,16'h00ae,16'h006a,-16'h0098,-16'h016a,-16'h005f,16'h00ea,-16'h0082,-16'h007d,16'h0099,-16'h016a,-16'h0009,16'h01b0,-16'h0029,-16'h0042,16'h0087,16'h00ae,16'h00b5,-16'h0080,16'h013a,-16'h0042,16'h00d4,-16'h0037,16'h017b,-16'h01b1,-16'h0066,-16'h01a5,16'h0039,16'h0006,16'h013a,-16'h00e6,-16'h000a,-16'h001d,16'h0027,16'h0175,16'h0140,-16'h0387,16'h00e4,16'h012f,16'h009d,16'h00c7,16'h000a,16'h0171,16'h0140,16'h008a,16'h0103,-16'h0023,16'h0138,16'h0003,16'h0046,16'h00aa,-16'h00e5,-16'h0020,-16'h0063,16'h0063,16'h00e9,16'h01bd,16'h0063,-16'h01b7,16'h0090,-16'h00ab,-16'h0190,-16'h0008,16'h01a5,16'h016b,16'h00c2,16'h0069,-16'h013b,16'h0039,-16'h0016,16'h00d6,16'h0024,-16'h0059,16'h00d8,-16'h01f8,-16'h0065,16'h0177,16'h003b,-16'h004d,16'h0097,-16'h0012,16'h0088,-16'h00bc,16'h007f,-16'h0058,16'h00c2,-16'h006e,16'h00f8,-16'h0178,16'h000d,-16'h023d,16'h005a,16'h0017,16'h0130,-16'h0082,-16'h00aa,16'h00b4,-16'h0059,16'h01aa,16'h00a7,-16'h02cc,16'h0134,16'h00ba,16'h00cc,16'h00f3,16'h00a2,16'h00f2,16'h0163,16'h00ef,16'h00d7,-16'h00e9,16'h00d7,16'h003a,-16'h009b,16'h00bd,-16'h009c,16'h001d,-16'h004c,16'h011a,16'h00e9,16'h0254,-16'h0208,-16'h0141,-16'h005a,16'h0004,-16'h0021,16'h0074,16'h0095,16'h011b,16'h00c1,16'h00f2,-16'h00c6,16'h013e,16'h0059,-16'h0116,16'h0076,-16'h0033,16'h00db,-16'h0135,-16'h0049,16'h01a6,16'h0081,-16'h0006,16'h0072,-16'h001c,16'h000c,-16'h0073,16'h00bd,16'h0013,16'h00e1,-16'h014f,16'h004c,-16'h0005,-16'h0020,-16'h01f7,16'h00a3,16'h00da,16'h0177,-16'h00f2,16'h0002,16'h00a7,-16'h00a1,16'h01cc,16'h009d,-16'h0239,16'h012b,16'h00df,16'h00ab,16'h002f,16'h0000,16'h0111,16'h00a7,16'h010f,16'h0109,-16'h00e5,16'h00d5,16'h0048,-16'h0120,16'h00ca,-16'h007a,16'h0037,-16'h0043,16'h0149,16'h0017,16'h024b,-16'h01ff,-16'h0132,-16'h0004,-16'h0033,16'h013b,16'h00e4,-16'h00e0,16'h001b,16'h00d3,16'h006a,16'h0027,16'h009a,16'h008e,-16'h0232,-16'h0054,16'h0045,16'h0105,-16'h00f2,-16'h0057,16'h0133,16'h00d4,16'h000e,16'h0071,16'h0010,16'h0023,-16'h0082,16'h013b,-16'h0042,16'h00cb,-16'h00d2,-16'h0030,16'h0098,16'h009a,-16'h007b,16'h00a3,16'h00de,16'h00d7,-16'h0089,-16'h0015,16'h0015,-16'h0038,16'h0032,16'h0092,-16'h0212,16'h011d,16'h0072,-16'h0018,16'h0034,16'h0033,16'h00d8,16'h00a6,16'h012e,16'h0190,-16'h00aa,16'h0075,16'h006a,-16'h0080,16'h014e,-16'h0030,16'h0047,16'h0006,16'h00bd,-16'h0050,16'h01c7,-16'h0200,-16'h018b,16'h000f,-16'h007a,16'h01c8,16'h009e,-16'h016e,-16'h01f8,16'h0112,16'h0052,16'h0132,16'h0014,-16'h001d,-16'h01f7,-16'h0074,-16'h0046,16'h00a8,-16'h004e,-16'h0020,16'h00cd,16'h00e4,-16'h0015,16'h0109,16'h001f,-16'h0017,-16'h00ca,16'h01bf,-16'h004c,16'h0062,-16'h00ac,16'h0035,16'h01cd,16'h0060,-16'h0041,16'h0113,16'h004d,16'h0027,-16'h0090,-16'h005b,16'h00b1,-16'h0027,-16'h0032,16'h007c,-16'h01cc,16'h013a,16'h0069,-16'h004f,16'h0079,16'h003d,16'h012f,16'h0000,16'h00dc,16'h00bf,-16'h001e,16'h0027,-16'h003e,16'h007d,16'h016c,16'h0040,16'h002d,16'h00c7,16'h0053,-16'h0047,16'h0248,-16'h013f,-16'h0200,-16'h003f,-16'h0102,16'h01b8,16'h0032,-16'h0168,-16'h0210,16'h00da,16'h000f,16'h009a,-16'h004b,-16'h0013,-16'h00ed,-16'h0009,-16'h0070,16'h001e,16'h007d,-16'h000d,16'h0089,16'h00b7,16'h0087,16'h00d3,16'h007c,-16'h008c,-16'h0010,16'h01a5,-16'h006a,-16'h0027,-16'h00c5,-16'h0044,16'h01fe,-16'h0021,-16'h0051,16'h0109,16'h0029,16'h0043,-16'h00b3,-16'h005e,16'h0046,-16'h0066,16'h002c,16'h0048,-16'h019d,16'h00a3,16'h0055,-16'h00c9,16'h00cc,-16'h003f,16'h00fc,16'h006d,16'h00f7,16'h00fe,-16'h0010,-16'h0031,-16'h001a,16'h0005,16'h0135,16'h001b,16'h006b,16'h0097,-16'h0061,-16'h0058,16'h01ae,-16'h00de,-16'h01ce,-16'h002b,-16'h00a6,16'h00d9,-16'h0077,-16'h017e,-16'h0289,16'h00d5,16'h0080,16'h0083,16'h00a3,-16'h006f,16'h005f,-16'h0058,16'h00a3,16'h00c5,-16'h0001,16'h0036,16'h0022,16'h0069,16'h0033,16'h012f,16'h0007,16'h0019,-16'h0038,16'h018d,-16'h001c,16'h003c,-16'h0166,-16'h0005,16'h019e,-16'h0029,16'h0014,16'h0099,16'h007c,16'h001b,16'h0013,-16'h0090,16'h008e,-16'h004d,16'h00a8,16'h0064,-16'h0142,16'h00ab,16'h007d,-16'h0163,16'h003e,-16'h0139,16'h017e,16'h0075,16'h012d,16'h0187,-16'h001f,-16'h004e,16'h0090,-16'h0032,16'h017c,16'h004d,16'h00c6,16'h00b9,-16'h0062,16'h001c,16'h019e,16'h0077,-16'h01b4,16'h0111,-16'h007c,16'h0072,-16'h0026,-16'h00c3,-16'h019c,16'h00d7,16'h010b,16'h001b,16'h014c,-16'h009b,16'h014d,-16'h008e,16'h00af,16'h00b0,-16'h0058,-16'h0030,16'h002e,16'h012f,16'h000d,16'h013e,16'h005d,16'h008c,-16'h0026,16'h016a,16'h003d,16'h0075,-16'h00d0,-16'h00ae,-16'h012e,-16'h007b,16'h0076,16'h00bf,16'h0089,16'h003a,-16'h0099,-16'h0101,16'h005c,16'h0056,16'h0180,16'h009c,-16'h01b8,16'h0079,16'h0022,-16'h011e,-16'h0045,-16'h0250,16'h008a,16'h00de,16'h00b5,16'h0190,-16'h0074,-16'h0072,16'h0001,-16'h00a6,16'h0132,-16'h0026,16'h0054,16'h00e4,-16'h0055,-16'h0034,16'h013b,16'h00ad,-16'h0107,16'h00e9,-16'h0004,-16'h0058,-16'h00b5,-16'h0036,-16'h0113,16'h0127,16'h00be,-16'h011b,16'h00a2,-16'h0084,16'h00c7,-16'h0076,16'h007d,16'h0092,-16'h00a0,16'h003d,-16'h003c,16'h0166,-16'h000d,16'h00e9,16'h005b,16'h00de,-16'h009d,16'h019f,-16'h001c,16'h0073,-16'h0050,-16'h0146,-16'h0221,-16'h00a8,16'h0114,16'h0066,16'h0112,16'h002c,-16'h006b,-16'h007d,16'h007c,16'h00cb,16'h020a,16'h0031,-16'h0209,-16'h0002,16'h006b,-16'h0112,-16'h008c,-16'h034f,16'h00a5,16'h008a,16'h0022,16'h0123,-16'h0050,-16'h002a,-16'h0015,-16'h0064,16'h0181,16'h0033,16'h004e,16'h009b,-16'h007b,16'h006a,16'h0135,16'h0042,16'h000b,16'h013e,16'h0058,-16'h00cc,-16'h00d7,-16'h0020,-16'h006f,16'h0155,16'h00b8,-16'h012c,-16'h000d,-16'h00e0,16'h007b,-16'h005c,16'h00bc,16'h0084,-16'h005c,16'h008d,-16'h0046,16'h00da,-16'h0017,16'h0064,16'h0107,16'h00da,-16'h00a9,16'h0188,-16'h0053,16'h0147,16'h0012,-16'h00e8,-16'h02aa,-16'h0051,16'h010a,-16'h003c,16'h00b3,16'h00c5,-16'h00a1,-16'h0048,16'h00c1,16'h0014,16'h01fd,16'h009f,-16'h0186,-16'h000d,16'h0087,-16'h00db,16'h0041,-16'h04ac,16'h0066,16'h00de,16'h0051,16'h016e,-16'h00c2,-16'h003f,16'h000f,16'h0034,16'h013e,16'h0032,16'h0099,16'h006f,-16'h0023,16'h00e4,16'h00f5,16'h00fb,-16'h00f4,16'h01b6,16'h0041,16'h0048,16'h0019,-16'h012b,16'h0079,16'h010d,16'h0061,-16'h010a,-16'h0033,-16'h00c6,16'h0005,16'h0028,16'h0196,16'h012b,16'h0131,16'h0079,16'h003d,16'h0035,-16'h010d,16'h00e1,16'h0058,16'h0144,-16'h0004,16'h01a9,-16'h00d2,16'h008b,16'h0008,-16'h014b,-16'h0178,-16'h0042,16'h00d0,-16'h0055,16'h018a,16'h011f,-16'h00b1,-16'h006c,16'h0170,16'h005e,16'h0200,16'h0087,-16'h019f,16'h001a,16'h00f0,-16'h0111,16'h0060,-16'h05e1,16'h002d,16'h0043,16'h0057,16'h0142,-16'h003d,16'h000a,-16'h0069,-16'h000b,16'h0137,-16'h0045,16'h0018,16'h00a3,-16'h000a,16'h00c9,16'h011c,16'h00ff,-16'h004d,16'h018c,16'h00ad,16'h0040,16'h00c9,-16'h00e4,16'h0047,16'h0154,16'h001a,-16'h0020,-16'h0141,-16'h0024,-16'h0055,-16'h0072,16'h0087,16'h0074,16'h0177,16'h00d8,16'h00de,-16'h001d,-16'h00b7,16'h0193,16'h006d,16'h0106,-16'h006c,16'h011f,-16'h0076,16'h0142,-16'h0016,-16'h019c,16'h0061,-16'h00ab,16'h00ac,-16'h008c,16'h0154,16'h00f6,-16'h0185,-16'h008a,16'h00d6,16'h0012,16'h0141,16'h00d6,-16'h010a,16'h00df,16'h00e6,-16'h00c4,16'h0167,-16'h07cb,16'h0092,16'h0038,16'h0071,16'h0143,-16'h0085,16'h0030,-16'h002a,16'h0024,16'h00f2,-16'h000b,-16'h005d,-16'h0026,-16'h0027,16'h0029,16'h0100,16'h00a0,-16'h006a,16'h0091,16'h00c3,16'h0076,16'h015b,-16'h00eb,16'h0033,16'h0172,-16'h0040,16'h0062,-16'h0094,16'h0058,-16'h00f2,-16'h0094,16'h008d,16'h0082,16'h010f,16'h00b2,16'h00c1,16'h0060,-16'h0171,16'h0165,16'h0042,16'h00b7,-16'h0073,16'h0101,-16'h00a1,16'h00e3,-16'h0056,-16'h014d,16'h0164,-16'h0055,16'h00fc,-16'h0025,16'h00de,16'h0125,-16'h01bb,16'h0063,16'h00b3,16'h0097,16'h00f6,16'h007d,-16'h0119,16'h00ca,16'h00b0,-16'h00b1,16'h00e4,-16'h07d1,16'h003d,-16'h003e,-16'h0046,16'h0166,-16'h0079,16'h00e8,16'h00b8,16'h00a2,16'h00d6,16'h005a,-16'h0010,16'h015d,16'h0044,-16'h0047,16'h00e6,16'h0086,-16'h0015,-16'h02df,16'h011c,-16'h0014,16'h0164,-16'h007e,16'h0083,16'h018e,-16'h0029,16'h0153,-16'h00f8,16'h0004,-16'h00eb,-16'h00ea,16'h001a,16'h0042,16'h005a,16'h011b,16'h0110,16'h006f,-16'h02c0,16'h011d,-16'h002a,16'h0095,-16'h00bf,16'h00f8,16'h0037,16'h001f,-16'h0061,-16'h00f1,16'h00df,-16'h0007,16'h00c3,-16'h0045,16'h0065,16'h0094,-16'h01b2,-16'h000a,16'h0033,-16'h0013,16'h0004,-16'h006e,-16'h010b,16'h0176,16'h0025,-16'h0043,16'h0096,-16'h070c,16'h006b,16'h005f,16'h006b,16'h010f,16'h0025,16'h00c3,16'h003a,16'h0071,16'h0091,16'h009a,16'h0052,16'h0046,-16'h0007,-16'h012a,16'h011c,16'h0040,-16'h005c,-16'h08c0,16'h012b,16'h000a,16'h01ca,-16'h013e,16'h0069,16'h017d,16'h0021,16'h019e,-16'h0086,16'h007c,-16'h00a6,-16'h00e3,16'h0038,16'h0006,-16'h0003,16'h00d8,16'h0097,16'h00eb,-16'h03b1,16'h0133,-16'h00c5,16'h006a,-16'h00bd,16'h014a,16'h002a,-16'h0096,-16'h00bd,-16'h00ab,16'h0051,16'h0046,16'h0061,-16'h00ba,-16'h01f7,16'h001f,-16'h015c,-16'h003a,16'h0059,-16'h006e,16'h00c5,-16'h0055,-16'h00bc,16'h01a9,16'h0044,-16'h003a,16'h00a6,-16'h0531,16'h0029,16'h004d,16'h0074,16'h006e,16'h009c,16'h001f,16'h00bf,16'h0020,16'h0113,16'h0029,16'h00ce,-16'h01dc,-16'h009d,-16'h023b,16'h0173,-16'h007f,-16'h010f,-16'h0a70,16'h0171,16'h009e,16'h0221,-16'h0176,-16'h0042,16'h00f3,16'h015b,16'h01d8,-16'h00ec,16'h0014,-16'h0047,-16'h0158,16'h005f,16'h0081,16'h004b,16'h00dc,-16'h002f,16'h0023,-16'h0300,16'h00a7,-16'h00b3,16'h00d1,-16'h00d8,16'h0191,16'h0058,16'h0023,-16'h00b2,16'h0008,-16'h0087,16'h009b,16'h019b,-16'h003a,-16'h0760,16'h0084,-16'h01c7,-16'h0060,16'h009b,-16'h013d,16'h014c,16'h0025,-16'h0078,16'h0156,-16'h0059,16'h001a,16'h0084,-16'h0425,16'h00e0,16'h00c0,16'h007d,16'h0050,16'h00b9,-16'h004d,16'h001e,-16'h002e,16'h0133,16'h00d3,16'h001d,-16'h02cd,-16'h0068,-16'h033a,16'h00b5,-16'h00e4,-16'h00ec,-16'h0539,16'h0170,16'h00d8,16'h00f3,-16'h01e5,-16'h00cb,16'h0121,16'h0098,16'h0124,16'h0001,16'h000b,16'h00d7,-16'h00d6,16'h0047,16'h008b,16'h0084,16'h0126,16'h0037,16'h0015,-16'h0308,16'h00c4,-16'h00f8,16'h005e,16'h0027,16'h014f,16'h000c,16'h0086,16'h003d,16'h0037,-16'h0077,16'h001f,16'h00f9,-16'h00b9,-16'h0886,16'h0063,-16'h0137,16'h000b,16'h0010,-16'h01c1,16'h0175,16'h0030,-16'h005e,16'h0154,-16'h003d,-16'h0056,16'h006b,-16'h02fc,16'h005c,16'h0194,16'h003d,16'h003d,16'h0119,-16'h0089,-16'h0054,-16'h000f,16'h00b8,-16'h000f,-16'h0008,-16'h021e,-16'h0092,-16'h03f5,16'h012d,-16'h0113,-16'h009e,-16'h02ef,16'h0185,16'h001e,-16'h0340,-16'h0165,-16'h018d,16'h0140,-16'h005b,16'h019e,16'h00a3,-16'h0025,16'h0117,-16'h00d9,16'h00f6,16'h0054,16'h0019,16'h01ae,-16'h000c,16'h005d,-16'h033e,16'h003d,-16'h0111,-16'h005a,16'h00f2,16'h010f,16'h0066,16'h0095,16'h0111,16'h0042,16'h0051,16'h0011,16'h00ee,16'h0001,-16'h0498,16'h00f2,-16'h012b,-16'h00aa,16'h005b,-16'h016a,16'h0161,16'h0043,-16'h0018,16'h00e6,-16'h0068,-16'h0100,-16'h00e7,-16'h02ac,16'h00d1,16'h0257,16'h00b5,-16'h0043,16'h009c,-16'h004f,-16'h009b,16'h0050,16'h0121,-16'h0060,16'h0006,-16'h01ee,-16'h0012,-16'h0340,16'h00e6,-16'h0058,-16'h00ea,-16'h0165,16'h01af,16'h005d,-16'h065a,-16'h00e9,-16'h02b0,16'h0050,-16'h0012,16'h01cc,16'h0045,16'h002b,16'h00b4,-16'h0115,16'h00a3,-16'h0006,-16'h0004,16'h0210,-16'h0018,-16'h000a,-16'h02e4,16'h000f,-16'h0122,-16'h001e,16'h0242,16'h00f3,16'h014a,16'h00dd,16'h01ee,-16'h0061,-16'h0030,-16'h009c,16'h00c4,16'h0012,-16'h01e8,16'h010e,-16'h01bb,-16'h00e0,16'h0062,-16'h008f,16'h0189,16'h009f,-16'h0010,-16'h0076,-16'h0077,-16'h00b8,-16'h011b,-16'h0227,16'h005d,16'h0278,16'h0050,-16'h016e,16'h0147,-16'h000d,-16'h0136,16'h0075,16'h019b,-16'h0067,16'h0080,-16'h013e,-16'h00bc,-16'h020f,16'h00b2,-16'h0053,-16'h00d6,-16'h0026,16'h0216,16'h0081,-16'h062d,-16'h0031,-16'h027d,16'h0063,-16'h0100,16'h00eb,16'h0088,16'h0042,16'h0074,-16'h0031,16'h00b0,-16'h0007,16'h0007,16'h010e,16'h00cd,16'h0098,-16'h0232,-16'h00c8,-16'h0027,-16'h000e,16'h0258,16'h00ff,16'h016d,16'h00c9,16'h0272,16'h0039,-16'h0019,-16'h0036,16'h00e5,-16'h0013,-16'h00a3,-16'h005b,-16'h00cf,-16'h0043,16'h000c,-16'h002c,16'h017c,-16'h0001,-16'h000d,-16'h01d4,-16'h00cc,-16'h000c,-16'h0132,-16'h0273,-16'h0087,16'h021a,16'h0081,-16'h003e,16'h0087,16'h00cd,-16'h01b1,16'h0125,16'h01b7,-16'h0069,16'h00a8,-16'h00e0,-16'h0085,-16'h0133,16'h00c0,-16'h0074,-16'h00c3,16'h009e,16'h01ea,16'h00d9,-16'h03a9,-16'h0048,-16'h023e,16'h009f,-16'h012a,-16'h0025,16'h000c,16'h00c4,16'h0049,16'h0014,16'h0089,16'h000c,16'h016c,16'h00ff,16'h0170,16'h0045,-16'h0240,-16'h0034,-16'h0092,-16'h0071,16'h0135,16'h0162,16'h0065,16'h0003,16'h01fb,16'h0017,-16'h004e,-16'h008d,16'h0074,16'h0052,16'h0010,-16'h0132,-16'h00fe,16'h00cf,16'h012a,16'h0095,16'h00bb,16'h00cf,-16'h0138,16'h0086,16'h0106,16'h0045,16'h00f9,16'h017a,-16'h0071,16'h025f,-16'h00c6,16'h0249,-16'h0025,-16'h0012,16'h0097,16'h0021,16'h002a,16'h0026,-16'h015c,-16'h012f,16'h0036,16'h01ef,-16'h00bc,-16'h00aa,-16'h0210,16'h0059,-16'h0055,16'h0084,-16'h0021,16'h030f,16'h018f,16'h0129,16'h009e,-16'h0152,-16'h006c,16'h0179,-16'h0054,-16'h005f,16'h01d6,16'h001f,16'h004e,16'h007d,16'h0025,16'h0054,-16'h001a,16'h002d,16'h00e6,16'h0093,-16'h0060,16'h01fe,-16'h0043,16'h0050,16'h00b6,-16'h008f,16'h0057,-16'h00a9,-16'h0111,-16'h00f6,-16'h0085,16'h0201,-16'h003f,16'h0132,16'h00e1,16'h00d7,16'h00d9,16'h008c,-16'h0186,16'h00df,16'h00c0,16'h0061,16'h010e,16'h012b,16'h0004,16'h0263,-16'h014b,16'h01e9,-16'h0010,16'h0018,16'h0096,16'h009c,-16'h003c,16'h0032,-16'h0165,-16'h0094,16'h0034,16'h00fa,16'h0033,-16'h0016,-16'h02fd,16'h002e,16'h002a,16'h00ae,-16'h00bc,16'h0371,16'h01d2,16'h0062,16'h0021,-16'h0109,-16'h0085,16'h00f1,-16'h005b,-16'h006b,16'h020e,-16'h0022,16'h0028,16'h0077,16'h008c,-16'h002f,16'h002e,-16'h001d,16'h0014,16'h0080,-16'h0095,16'h015f,16'h0003,16'h0078,16'h0120,16'h0091,16'h0165,-16'h003c,-16'h015b,-16'h016b,-16'h00d3,16'h0123,16'h001b,16'h0105,16'h010a,16'h00c6,16'h00cc,16'h00d2,-16'h01ec,16'h011c,16'h00ba,-16'h0023,16'h0068,16'h00a6,16'h015f,16'h0280,-16'h023b,16'h017b,-16'h0008,16'h0081,-16'h000a,16'h00e3,-16'h0083,-16'h007e,-16'h0137,-16'h00b8,16'h0027,16'h0039,-16'h0051,-16'h0001,-16'h03ac,-16'h006a,-16'h009b,-16'h0002,-16'h003d,16'h0300,16'h0234,16'h0101,-16'h0016,-16'h0158,-16'h004c,-16'h0083,-16'h00fb,-16'h002e,16'h0259,-16'h007e,-16'h00d1,16'h0016,16'h00fd,-16'h0018,16'h005c,16'h00b6,16'h0029,16'h0073,-16'h00eb,16'h00c7,-16'h0001,16'h0013,16'h020f,16'h0154,16'h01d3,16'h001e,-16'h0110,-16'h017e,-16'h0004,16'h0040,-16'h003c,16'h00f2,16'h00cb,16'h00a0,16'h0146,16'h00b8,-16'h01ca,16'h0157,16'h0115,-16'h0009,16'h000f,16'h0063,16'h01f2,16'h0196,-16'h0159,-16'h0004,16'h001c,16'h005e,-16'h0083,16'h0021,-16'h0109,-16'h00d6,-16'h00af,-16'h0044,-16'h0111,-16'h0001,16'h00c7,16'h00b1,-16'h0328,-16'h0003,-16'h00e6,-16'h0004,-16'h00cc,16'h0266,16'h0154,16'h0032,-16'h00ab,-16'h0021,-16'h0001,-16'h00fa,-16'h009f,-16'h005f,16'h01ff,-16'h00da,-16'h0025,16'h008d,16'h00c0,-16'h0025,16'h0013,16'h0069,16'h0066,16'h00a5,-16'h00f4,16'h005d,16'h0016,-16'h007e,16'h0189,16'h01d1,16'h0117,-16'h001c,-16'h009c,-16'h0145,16'h0007,16'h0007,-16'h00c5,16'h01c2,16'h0032,16'h0128,16'h0166,16'h0127,-16'h01f6,16'h0200,16'h0090,16'h001a,16'h001e,16'h001b,16'h01e9,16'h0116,-16'h0107,-16'h00e2,16'h0020,16'h0018,-16'h00a4,16'h005b,-16'h019a,-16'h0017,-16'h004c,16'h0020,-16'h01f9,-16'h000d,16'h01a1,16'h012b,-16'h01a5,16'h00ab,-16'h013f,16'h009e,-16'h000a,16'h0172,16'h0103,16'h0013,-16'h00b9,16'h003f,16'h000d,-16'h0115,-16'h00b1,-16'h00c9,16'h0227,-16'h013f,16'h0028,16'h0063,16'h0084,-16'h0026,16'h002a,16'h006a,16'h006a,16'h00a5,-16'h01a6,16'h005b,-16'h0073,-16'h0031,16'h01ae,16'h0180,16'h0054,-16'h00d0,-16'h0151,-16'h0142,16'h005a,16'h00e9,-16'h0118,16'h017f,-16'h0021,16'h00b5,16'h0179,16'h016e,-16'h0188,16'h0225,16'h011c,16'h00b5,-16'h0025,-16'h0005,16'h0235,16'h00cb,-16'h0138,-16'h0150,16'h0053,-16'h0084,-16'h00ae,16'h0019,-16'h01e1,-16'h006b,-16'h0062,16'h009a,-16'h01be,-16'h005d,16'h01c8,16'h0205,-16'h0013,16'h0033,-16'h012e,-16'h0055,16'h003f,16'h01c2,16'h00e2,16'h00bd,-16'h00d9,16'h0120,-16'h008d,-16'h0203,-16'h00de,-16'h009d,16'h0219,-16'h00ea,-16'h0046,16'h0036,16'h0124,-16'h0022,16'h0000,16'h00d3,16'h0008,-16'h0006,-16'h008c,16'h0078,-16'h0052,-16'h007a,16'h010b,16'h0209,-16'h0028,-16'h010b,-16'h018c,-16'h00f0,-16'h001b,16'h00a5,-16'h014b,16'h0172,16'h001e,16'h0048,16'h014e,16'h0143,-16'h017a,16'h0238,16'h00f5,16'h00c0,16'h005e,-16'h001a,16'h0207,16'h00e4,-16'h00fe,-16'h00e3,16'h0079,-16'h00b3,16'h001a,16'h0072,-16'h0174,-16'h0082,-16'h0059,16'h0102,-16'h00e5,16'h008a,16'h01fd,16'h015d,-16'h0111,16'h0087,-16'h0138,-16'h00cf,16'h00d1,16'h01b4,16'h00b9,16'h0097,-16'h002b,16'h00b7,-16'h0190,-16'h0118,16'h00d1,-16'h009f,16'h0142,-16'h0077,-16'h0090,16'h0005,16'h00fa,16'h0013,-16'h0027,16'h00ae,-16'h0024,16'h0065,-16'h0043,16'h0089,-16'h00ba,-16'h009b,16'h007c,16'h0104,-16'h013e,-16'h00fa,-16'h013f,-16'h0099,16'h0001,16'h011f,-16'h0110,16'h0109,-16'h0060,16'h004b,16'h0169,16'h0069,-16'h01a0,16'h023d,16'h012c,16'h0126,16'h0071,16'h0034,16'h024f,16'h00ad,16'h0011,-16'h00c2,16'h0060,16'h000f,16'h0063,16'h013d,-16'h007c,-16'h010e,-16'h0039,16'h011b,16'h0008,16'h0098,16'h022f,16'h012c,-16'h014f,-16'h0020,-16'h0100,-16'h011c,16'h0099,16'h0141,16'h00a5,16'h00cb,16'h00b4,-16'h00ce,-16'h0128,-16'h0089,16'h00f9,-16'h005d,16'h014a,16'h0030,-16'h013b,-16'h0025,16'h00f5,16'h0015,-16'h0046,16'h00a3,16'h005b,16'h00c2,16'h002d,16'h0071,-16'h00a7,16'h0018,16'h0021,16'h00b0,-16'h0145,-16'h001f,-16'h01cf,-16'h002c,-16'h000d,16'h012c,-16'h0154,16'h0062,-16'h0084,16'h000f,16'h0147,-16'h002a,-16'h0193,16'h01aa,16'h0153,16'h0075,16'h006d,16'h0054,16'h021f,16'h00e9,16'h00f0,-16'h00f4,-16'h0016,16'h007e,16'h0064,16'h00ee,16'h003b,-16'h00ed,16'h0032,16'h0030,-16'h0005,16'h007f,16'h01be,16'h0035,-16'h018c,16'h0045,-16'h00dd,-16'h01b8,16'h0013,16'h01cf,16'h00c3,16'h0089,16'h0149,-16'h01be,16'h0011,16'h006a,16'h00aa,16'h001d,16'h00ad,16'h0017,-16'h0136,-16'h006e,16'h00e7,16'h00a4,-16'h0079,16'h0066,-16'h0048,16'h0079,16'h003a,-16'h0073,-16'h0089,16'h0077,-16'h008e,16'h0059,-16'h00c0,16'h0041,-16'h0265,16'h003d,16'h005b,16'h0107,-16'h00a1,16'h003e,-16'h0011,-16'h007c,16'h01a9,-16'h00f6,-16'h01f9,16'h01f7,16'h0097,16'h0012,16'h008b,-16'h0056,16'h01db,16'h005f,16'h0147,-16'h0045,-16'h00ca,16'h00ae,16'h00a0,-16'h000c,16'h00ac,-16'h0109,16'h0048,-16'h0099,16'h0016,16'h001e,16'h023c,-16'h015f,-16'h00e0,16'h0002,-16'h010e,-16'h00be,16'h00d3,16'h017d,16'h00c8,16'h00b1,16'h0042,-16'h00b2,16'h005f,16'h00e1,-16'h013d,16'h0000,16'h009f,-16'h002d,-16'h013d,-16'h013b,16'h00d9,-16'h0040,-16'h0033,16'h002b,16'h0032,16'h0091,-16'h0022,-16'h000a,-16'h0097,16'h00f3,-16'h010b,-16'h001a,-16'h0042,16'h0065,-16'h01df,16'h008e,16'h00c8,16'h0134,-16'h00dd,16'h0046,-16'h0074,-16'h0050,16'h0192,-16'h00af,-16'h012e,16'h02a3,16'h00be,16'h002d,16'h007b,-16'h0093,16'h0247,16'h009d,16'h00f6,-16'h0016,-16'h00fe,16'h00d7,16'h003c,16'h0047,16'h00f0,16'h0000,-16'h002a,-16'h0039,16'h002c,16'h0012,16'h020f,-16'h016b,-16'h008c,-16'h0032,-16'h012a,16'h00a5,16'h0129,16'h0124,-16'h00c6,16'h00b5,16'h00cf,16'h0040,16'h007d,16'h0072,-16'h02aa,-16'h0023,16'h00be,16'h005e,-16'h0118,-16'h00c6,16'h006d,16'h0094,16'h0010,16'h0111,16'h0012,16'h0086,-16'h0078,16'h0032,-16'h003d,16'h013d,-16'h00dd,-16'h004f,16'h00bc,16'h007e,-16'h01d7,16'h0065,16'h0125,16'h00b6,-16'h0105,16'h0014,-16'h0113,-16'h0069,16'h0116,16'h0034,-16'h01f9,16'h0293,16'h003f,-16'h0095,16'h0060,-16'h0183,16'h022c,16'h0087,16'h0147,-16'h002f,-16'h00b0,16'h0093,16'h0058,16'h0096,16'h0147,-16'h002c,-16'h000b,16'h001b,16'h0095,16'h0033,16'h024d,-16'h00fe,-16'h0056,-16'h0036,-16'h0162,16'h018f,16'h005d,16'h00b5,-16'h01dc,16'h011f,16'h0059,16'h00cc,-16'h00b8,16'h0001,-16'h0222,-16'h00d2,16'h00db,-16'h0050,-16'h0026,-16'h00b2,-16'h0025,16'h0097,-16'h00a8,16'h00ff,16'h0009,16'h0083,-16'h00c7,16'h00cf,-16'h00a7,16'h004a,-16'h0012,16'h0013,16'h010a,16'h0089,-16'h0205,16'h0048,16'h0121,16'h00a6,-16'h0105,-16'h004b,-16'h00b3,16'h0060,16'h004c,16'h0030,-16'h01ac,16'h02d4,16'h0002,-16'h00df,16'h00b8,-16'h025a,16'h01be,16'h002d,16'h0125,-16'h00b2,-16'h0028,16'h007b,16'h002b,16'h010a,16'h0162,-16'h0008,-16'h002b,16'h004b,-16'h001e,16'h0028,16'h0249,-16'h0135,-16'h018f,-16'h0013,-16'h01bb,16'h0160,-16'h000c,16'h00a3,-16'h0236,16'h0146,-16'h000a,16'h008a,-16'h0072,-16'h005c,-16'h014a,-16'h00b5,16'h00ad,-16'h000d,16'h0033,-16'h00ff,16'h000d,16'h00b6,-16'h0033,16'h00df,-16'h0017,16'h0036,-16'h00b0,16'h0120,-16'h00c1,16'h008a,-16'h0089,16'h0021,16'h0106,16'h005f,-16'h011c,-16'h0016,16'h015b,16'h000b,-16'h00ad,-16'h0083,-16'h009a,-16'h0022,16'h0047,-16'h0096,-16'h0109,16'h0273,16'h0002,-16'h017a,16'h00ff,-16'h02eb,16'h01f0,-16'h0014,16'h012a,-16'h00c4,-16'h0079,16'h0003,16'h0016,16'h00ea,16'h0120,-16'h002d,16'h006e,16'h008e,16'h003c,-16'h000a,16'h01aa,-16'h00d1,-16'h0243,16'h0004,-16'h0208,16'h0103,-16'h0045,16'h0003,-16'h0158,16'h00d9,-16'h0017,16'h0003,16'h0004,-16'h0129,-16'h0081,-16'h002c,16'h0008,-16'h0087,-16'h0013,-16'h0059,-16'h0005,16'h00f0,-16'h0063,16'h00f7,16'h0040,16'h006a,-16'h00a7,16'h00c5,-16'h011b,16'h008e,-16'h0078,-16'h005d,16'h00d6,-16'h0033,-16'h0055,16'h0009,16'h00e2,-16'h0033,-16'h00a8,-16'h00a8,-16'h0016,16'h0065,16'h0057,-16'h00ce,-16'h00d7,16'h018e,16'h004b,-16'h011c,16'h003d,-16'h0475,16'h01fb,16'h0010,16'h0163,-16'h00e7,-16'h00a3,-16'h0073,-16'h003e,16'h007b,16'h00b1,-16'h0003,16'h0071,16'h00b0,16'h0018,16'h0033,16'h0144,16'h000e,-16'h018a,16'h0089,-16'h02b1,16'h00e4,-16'h0013,-16'h0054,-16'h0115,16'h007b,16'h0024,-16'h00d4,16'h00a3,-16'h00f3,16'h00f5,-16'h003d,16'h005a,-16'h003c,-16'h00a9,-16'h005d,-16'h005b,16'h0100,-16'h0067,16'h00da,16'h0041,16'h00d3,-16'h00b7,16'h0166,-16'h00af,16'h0005,-16'h00e0,-16'h00f4,-16'h016d,-16'h0059,16'h0033,-16'h0018,16'h00b6,-16'h0044,-16'h00e1,-16'h0077,16'h003b,16'h00a4,16'h0106,-16'h011c,16'h0003,16'h0174,16'h004b,-16'h00d1,16'h0028,-16'h0574,16'h01ee,-16'h0018,16'h0135,-16'h0107,-16'h00e8,-16'h0094,-16'h0053,16'h0021,16'h0134,16'h0035,16'h00a7,16'h0085,16'h0018,16'h0083,16'h019c,16'h0006,-16'h004b,16'h011e,-16'h022a,16'h004f,-16'h0072,-16'h0065,-16'h0071,16'h00a2,16'h0053,-16'h012c,16'h0061,-16'h010c,16'h00bc,-16'h0108,16'h0086,-16'h0060,-16'h011c,-16'h0006,-16'h001b,16'h012e,-16'h0043,16'h00db,16'h007a,16'h00d8,-16'h0031,16'h0130,-16'h00b6,16'h0040,-16'h0067,-16'h0083,-16'h0286,-16'h00ef,16'h004a,16'h0011,16'h0130,-16'h003d,-16'h00dd,-16'h00a5,-16'h0036,16'h006e,16'h017c,-16'h00f2,-16'h0139,16'h0110,16'h0071,-16'h00af,-16'h0085,-16'h06f0,16'h01b7,-16'h0005,16'h00c9,-16'h00f5,-16'h00c6,-16'h009c,16'h0001,16'h0016,16'h00f9,16'h003b,16'h0002,16'h0057,-16'h006e,16'h0053,16'h01a2,16'h002b,-16'h0070,16'h017f,-16'h023d,-16'h010b,-16'h00d2,-16'h000e,-16'h0015,16'h011d,16'h00e3,-16'h01c2,16'h004a,-16'h0194,16'h00be,-16'h0011,16'h00a5,-16'h0021,-16'h0031,16'h009b,-16'h0019,16'h0106,-16'h0140,16'h0120,16'h006e,16'h0118,-16'h0067,16'h00f9,-16'h008c,16'h005e,-16'h00d0,-16'h0071,-16'h02b9,-16'h0190,16'h009b,-16'h0007,16'h0147,16'h000f,-16'h00af,-16'h007c,16'h0044,16'h0004,16'h019a,-16'h010d,-16'h00dc,16'h00ed,16'h00d8,-16'h0136,16'h000a,-16'h0787,16'h00f5,16'h0036,16'h003c,-16'h0119,-16'h00b7,-16'h006b,-16'h00b0,16'h007d,16'h0136,-16'h000c,16'h002c,16'h0039,-16'h009e,16'h00eb,16'h0140,16'h008d,-16'h013a,16'h015e,-16'h01e4,16'h0009,16'h0065,-16'h003c,-16'h0004,16'h00f4,16'h000d,-16'h00ed,-16'h0093,-16'h0133,-16'h0006,-16'h0026,16'h00f1,16'h0037,16'h00ff,16'h00e1,16'h0038,16'h0058,-16'h01fe,16'h0121,16'h003e,16'h0133,-16'h00a0,16'h00ab,-16'h00cd,16'h00c9,-16'h00df,-16'h014c,-16'h00fc,-16'h0137,16'h0117,-16'h0046,16'h00aa,16'h008f,-16'h010c,-16'h0062,-16'h0018,-16'h0020,16'h0194,16'h0060,-16'h0168,16'h00b4,16'h00ea,-16'h0090,16'h0065,-16'h08c3,16'h007b,-16'h004c,16'h005d,-16'h0081,-16'h0055,16'h0073,-16'h002d,16'h0023,16'h0155,16'h0052,16'h0002,16'h0064,-16'h0047,16'h00c1,16'h00f9,16'h010b,-16'h006f,16'h00b3,-16'h01be,16'h0053,16'h00d7,-16'h00ac,-16'h0007,16'h00d8,16'h0029,-16'h003e,-16'h00ce,-16'h00bd,-16'h0082,-16'h0042,16'h0190,16'h0011,16'h0169,16'h00ac,16'h0044,16'h0007,-16'h02c8,16'h00d8,-16'h001e,16'h005a,-16'h004f,16'h0043,-16'h0080,16'h0050,-16'h00cd,-16'h01ad,16'h0077,-16'h00c8,16'h00a7,-16'h0021,16'h0090,16'h0080,-16'h014c,-16'h00a2,16'h008e,-16'h0064,16'h0189,16'h00b5,-16'h013d,16'h010d,16'h00df,-16'h0068,16'h00f8,-16'h0894,16'h00b7,-16'h00f4,16'h00ab,-16'h0037,-16'h004a,-16'h002a,16'h001f,16'h0056,16'h018c,16'h007e,-16'h00d5,16'h0047,16'h0057,-16'h0063,16'h0119,16'h00c5,16'h0089,16'h0087,-16'h00f6,16'h0028,16'h0119,-16'h0193,16'h0077,16'h007c,16'h0026,16'h0077,-16'h0046,-16'h0050,-16'h013e,-16'h0082,16'h0109,16'h0041,16'h0149,16'h00d7,16'h0099,16'h0065,-16'h0304,16'h00e2,-16'h0047,16'h0084,-16'h003b,16'h0098,16'h0011,16'h0087,-16'h00a4,-16'h014e,16'h00bf,-16'h009e,16'h017b,16'h0017,-16'h0021,16'h00b5,-16'h00fc,16'h0015,16'h0093,16'h00b5,16'h00f8,16'h0005,-16'h020e,16'h01a3,16'h0135,16'h0025,16'h00b3,-16'h07a5,16'h0095,-16'h008c,-16'h0018,-16'h0045,16'h0004,16'h00ef,16'h0004,16'h0088,16'h011b,16'h00a3,-16'h0023,16'h006f,16'h0039,-16'h0109,16'h0106,16'h0076,16'h006f,-16'h02b4,-16'h00f7,-16'h009f,16'h0140,-16'h01d8,16'h005d,16'h007f,16'h0027,16'h0149,-16'h009b,16'h00e0,-16'h011f,-16'h002f,16'h0073,16'h000d,16'h0105,16'h0113,16'h0084,16'h0032,-16'h0472,16'h014c,-16'h0011,16'h0032,-16'h00c5,16'h00dc,-16'h000a,16'h001e,16'h0005,-16'h00d0,16'h014d,16'h0010,16'h0127,16'h0019,-16'h004b,16'h00b2,-16'h00eb,-16'h003b,16'h0017,-16'h0042,16'h00e8,-16'h0017,-16'h01e4,16'h0159,16'h0088,-16'h0063,16'h00e6,-16'h05ce,16'h0079,-16'h0064,16'h0038,-16'h0057,16'h002c,16'h0053,16'h001c,16'h00cb,16'h0161,16'h00b6,16'h0082,16'h0022,-16'h0031,-16'h0196,16'h015f,16'h003c,-16'h003b,-16'h0872,-16'h00a3,16'h0074,16'h0175,-16'h01f8,16'h0043,16'h00bd,16'h005f,16'h0168,-16'h0018,16'h00cf,-16'h0122,-16'h006f,16'h009b,-16'h0024,16'h0102,16'h018d,-16'h002f,16'h006a,-16'h03fc,16'h012c,-16'h00ae,16'h006d,-16'h013c,16'h00e0,16'h0032,-16'h0033,16'h0099,-16'h0008,-16'h0015,16'h00a9,16'h0165,16'h0000,-16'h02a5,16'h00dc,-16'h00be,-16'h00d9,16'h00c4,-16'h00a5,16'h0137,-16'h0062,-16'h0218,16'h011e,16'h008b,-16'h0037,16'h0092,-16'h042f,16'h0086,-16'h0032,-16'h0034,-16'h00c4,16'h00bb,16'h0040,16'h001b,16'h0087,16'h0192,16'h0074,16'h00bb,-16'h015b,-16'h0053,-16'h02ab,16'h017a,16'h005d,-16'h00d9,-16'h096f,-16'h00a7,16'h00bd,16'h01a3,-16'h0207,-16'h00d8,16'h00f7,16'h016e,16'h01c1,-16'h0080,16'h00fc,-16'h0016,-16'h008f,-16'h0005,16'h0054,16'h0072,16'h00e9,16'h0030,16'h002e,-16'h0304,16'h0072,-16'h0153,16'h0006,-16'h00b8,16'h018e,16'h00ec,-16'h002e,16'h0080,-16'h0017,-16'h008f,16'h00f9,16'h012f,-16'h004b,-16'h07a6,16'h0018,-16'h00ee,16'h00b5,16'h00a5,-16'h01d4,16'h0125,-16'h0034,-16'h01d9,16'h0112,16'h004d,-16'h0077,16'h0036,-16'h0337,16'h0111,16'h0028,16'h0004,-16'h008c,16'h00a8,16'h0046,-16'h000b,-16'h0047,16'h0137,16'h00db,-16'h0037,-16'h01ec,-16'h0006,-16'h03ab,16'h0171,16'h0014,-16'h010b,-16'h0544,16'h0022,16'h0130,16'h0053,-16'h01b7,-16'h00fa,16'h0114,16'h00eb,16'h014b,16'h0024,16'h00ae,16'h00ee,-16'h00f8,16'h007d,16'h007a,16'h0054,16'h0062,-16'h001d,-16'h001a,-16'h0280,16'h00a2,-16'h0182,-16'h0056,16'h0060,16'h0143,16'h00c2,-16'h0021,16'h0060,-16'h003a,-16'h00e6,16'h00ab,16'h01b4,16'h0039,-16'h06c8,16'h0066,-16'h00be,-16'h0044,16'h00c6,-16'h0201,16'h015a,16'h0029,-16'h011c,16'h0122,-16'h001f,-16'h0078,-16'h007f,-16'h02bb,16'h008a,16'h0114,16'h007a,-16'h00cd,16'h00ea,-16'h006e,-16'h0040,16'h002c,16'h0122,16'h001d,16'h0004,-16'h0202,-16'h0076,-16'h03b6,16'h0115,-16'h0033,-16'h011b,-16'h0299,16'h0034,16'h009a,-16'h02af,-16'h00d7,-16'h01db,16'h00bb,-16'h0036,16'h022c,16'h007e,16'h0053,16'h0141,-16'h003a,16'h00c3,16'h00a6,-16'h0025,16'h015f,-16'h002d,16'h0075,-16'h0276,16'h0011,-16'h0171,-16'h00d1,16'h015a,16'h00c8,16'h00cb,16'h003b,16'h011d,-16'h0056,-16'h0070,-16'h005b,16'h0187,-16'h000a,-16'h0395,16'h00c0,-16'h00ab,-16'h005f,16'h0057,-16'h016a,16'h0170,16'h006d,-16'h00b6,16'h00de,-16'h0057,-16'h0048,-16'h016b,-16'h0248,16'h0088,16'h01ff,16'h0000,-16'h012a,16'h00a6,-16'h001d,-16'h0133,16'h0099,16'h019e,-16'h0060,-16'h001a,-16'h019f,-16'h00c8,-16'h02ef,16'h0131,16'h0035,-16'h00d4,-16'h016b,16'h00e4,16'h00d7,-16'h05d1,-16'h00ec,-16'h0237,16'h0081,-16'h009b,16'h018e,16'h0018,16'h0075,16'h008c,-16'h00be,16'h0084,-16'h0022,16'h00df,16'h0120,16'h0096,16'h007b,-16'h0178,-16'h0031,-16'h012d,-16'h008c,16'h02d7,16'h016f,16'h014c,16'h002e,16'h0165,-16'h0063,-16'h00ce,-16'h00a4,16'h0118,16'h0077,-16'h01c5,16'h00a0,-16'h00b9,-16'h00ea,16'h001a,-16'h0092,16'h01bd,16'h007f,-16'h003b,-16'h002f,-16'h0062,-16'h0012,-16'h0180,-16'h01fa,-16'h006d,16'h0291,16'h0000,-16'h0172,16'h00fa,16'h000a,-16'h020b,16'h0182,16'h01b9,-16'h0096,16'h0045,-16'h01f2,-16'h0097,-16'h01d6,16'h0114,16'h0049,-16'h00f1,16'h0026,16'h0106,16'h00b0,-16'h051e,-16'h0083,-16'h01aa,16'h00dc,-16'h0166,16'h0123,16'h007c,16'h0013,16'h005c,-16'h002c,16'h00cb,-16'h0056,16'h00e6,16'h005f,16'h007e,16'h0000,-16'h019d,-16'h0049,-16'h006b,-16'h0079,16'h0286,16'h0183,16'h00d4,16'h00bb,16'h0283,16'h0065,-16'h0080,-16'h005e,16'h0104,-16'h0041,-16'h000e,-16'h0091,-16'h00f9,-16'h0014,16'h0039,-16'h003b,16'h0158,16'h0020,-16'h00f4,-16'h00f8,-16'h0021,16'h0068,-16'h0117,-16'h019b,-16'h008b,16'h02b8,16'h00e2,-16'h0004,16'h0031,16'h00cf,-16'h0143,16'h018d,16'h01b2,-16'h0023,16'h00a2,-16'h010c,-16'h0051,-16'h0156,16'h00e4,-16'h0064,-16'h0020,16'h008c,16'h0147,16'h011f,-16'h032b,-16'h000d,-16'h01be,16'h0093,-16'h0143,-16'h00ef,-16'h005f,16'h0078,16'h0073,16'h004c,16'h0115,16'h002a,16'h0282,16'h008c,16'h0104,16'h0067,-16'h014d,-16'h0001,-16'h0023,-16'h0075,16'h0125,16'h0178,-16'h006d,-16'h0023,16'h0180,16'h0035,-16'h00d0,-16'h006e,16'h0097,16'h0041,-16'h000f,-16'h017f,-16'h00cc,16'h0098,16'h0197,16'h009c,16'h004b,16'h002e,-16'h017b,16'h0150,16'h0119,-16'h0058,16'h0143,16'h0190,-16'h0009,16'h01d1,-16'h0120,16'h024a,-16'h0039,-16'h003b,16'h009c,16'h004a,-16'h0067,-16'h00c2,-16'h0181,-16'h00f2,16'h00b6,16'h0168,-16'h00ee,-16'h006e,-16'h0161,16'h00ed,-16'h004d,16'h00f5,-16'h009c,16'h026e,16'h012e,16'h0064,-16'h0002,-16'h0067,-16'h0037,16'h01da,-16'h00a0,16'h0052,16'h021c,16'h0065,16'h0056,16'h004a,16'h000b,16'h0084,16'h006e,16'h0011,16'h00bd,16'h017a,-16'h00a8,16'h01f5,16'h003e,16'h0074,16'h00f4,-16'h011d,-16'h0061,-16'h0157,-16'h011e,-16'h0142,-16'h008d,16'h0180,-16'h0003,16'h00da,16'h00c2,16'h007d,16'h00b7,16'h0053,-16'h016f,16'h0128,16'h0054,-16'h0051,16'h0100,16'h0195,16'h000f,16'h0226,-16'h011e,16'h01b6,-16'h0076,16'h0014,16'h006b,16'h0050,-16'h006d,-16'h00cb,-16'h0185,-16'h014d,16'h0041,16'h017b,-16'h009b,-16'h0061,-16'h0270,-16'h001b,-16'h001e,16'h009b,-16'h000e,16'h030c,16'h01e3,16'h00a3,16'h003d,-16'h006e,-16'h0082,16'h00d8,-16'h0046,-16'h002a,16'h01ff,-16'h0013,-16'h000d,-16'h0003,16'h003c,-16'h0029,16'h0053,16'h0008,16'h0075,16'h0065,-16'h007b,16'h0184,16'h0000,16'h0056,16'h0160,-16'h001e,16'h00d1,-16'h00ff,-16'h00d5,-16'h0161,-16'h009b,16'h01b4,16'h002b,16'h0072,16'h009b,16'h0043,16'h009b,-16'h002a,-16'h019d,16'h0209,16'h005b,-16'h0052,16'h007a,16'h00ae,16'h00ad,16'h02e2,-16'h017e,16'h00dd,-16'h0008,16'h00d8,-16'h0047,16'h00ab,-16'h0091,-16'h014a,-16'h011d,-16'h0099,-16'h002d,16'h002e,-16'h0072,16'h0016,-16'h02de,-16'h0018,-16'h0055,16'h00b0,-16'h0004,16'h0349,16'h0213,16'h00cd,-16'h0051,-16'h00d0,-16'h0031,16'h0083,-16'h0089,-16'h0032,16'h01d0,-16'h0027,16'h000d,-16'h0064,16'h007d,-16'h00df,16'h009e,16'h006a,16'h0042,16'h009b,-16'h0119,16'h006a,-16'h0043,16'h006f,16'h01c7,16'h0092,16'h01b0,-16'h0013,-16'h010b,-16'h00b2,-16'h0045,16'h00d4,-16'h0019,16'h00b1,16'h00d3,16'h0069,16'h00f3,-16'h0018,-16'h0170,16'h011b,16'h0126,-16'h0025,16'h0051,16'h003f,16'h0161,16'h023c,-16'h01f0,16'h0008,16'h0030,16'h001b,-16'h0023,16'h0073,-16'h00c5,-16'h00a2,-16'h0134,-16'h0003,-16'h0115,16'h008d,16'h005a,16'h006e,-16'h032d,16'h0064,-16'h00b2,16'h003d,-16'h0067,16'h026f,16'h016b,-16'h001c,-16'h00cf,-16'h0016,-16'h0052,-16'h0006,-16'h002c,-16'h0079,16'h0238,-16'h0135,-16'h005a,-16'h0055,16'h005c,-16'h005b,16'h0003,16'h0092,16'h000f,16'h007d,-16'h013f,16'h0099,-16'h005a,16'h0039,16'h0172,16'h0158,16'h00e9,-16'h0066,-16'h011e,-16'h00a7,16'h003f,16'h008e,-16'h0001,16'h010c,16'h00a4,16'h00bd,16'h0109,16'h0008,-16'h0086,16'h0188,16'h00c8,16'h0016,-16'h0016,-16'h0033,16'h015c,16'h0195,-16'h0128,-16'h0127,-16'h0028,-16'h001f,-16'h0021,16'h00ac,-16'h01e1,-16'h0099,-16'h00c5,16'h005a,-16'h018e,-16'h005c,16'h00dc,16'h00ef,-16'h0166,16'h0049,-16'h00e1,16'h002e,-16'h003c,16'h0154,16'h00d1,16'h0002,-16'h012c,16'h009d,-16'h0061,-16'h0128,-16'h0071,-16'h00de,16'h01e9,-16'h015f,16'h003a,-16'h0043,16'h007b,-16'h0082,16'h0025,16'h0134,-16'h00ea,16'h0027,-16'h0123,16'h0080,16'h0023,-16'h0031,16'h014a,16'h010d,16'h0044,-16'h0097,-16'h01a2,-16'h0099,16'h000d,16'h0045,-16'h000b,16'h013a,-16'h001d,16'h00ba,16'h0132,-16'h0083,-16'h0088,16'h01bf,16'h0121,16'h0001,16'h001c,-16'h00d0,16'h014f,16'h0179,-16'h0105,-16'h0242,16'h0013,16'h0000,-16'h001b,16'h008b,-16'h0227,-16'h004c,-16'h0051,16'h0100,-16'h019f,-16'h000b,16'h00f0,16'h0113,-16'h0043,16'h0019,-16'h00e9,16'h0019,16'h00fd,16'h017b,16'h00be,16'h0085,-16'h00ae,16'h008f,-16'h015a,-16'h01a0,16'h0006,-16'h0030,16'h0235,-16'h0150,-16'h005c,-16'h0095,16'h00d0,-16'h00b8,16'h0003,16'h0105,-16'h00dc,16'h006c,-16'h0137,16'h00d0,-16'h0011,16'h0052,16'h0173,16'h0174,-16'h0004,-16'h006c,-16'h026e,-16'h0054,16'h003c,16'h0134,-16'h0098,16'h00cb,-16'h0057,16'h0098,16'h0133,-16'h00ed,16'h0008,16'h01b7,16'h011d,16'h0016,-16'h004d,-16'h007a,16'h0194,16'h00a0,-16'h0093,-16'h02f6,16'h0072,-16'h001c,-16'h008e,16'h0058,-16'h021f,-16'h00a9,16'h0000,16'h0129,-16'h0140,16'h0046,16'h0198,16'h00d1,-16'h00af,-16'h0052,-16'h0094,-16'h0097,16'h00dc,16'h019c,16'h007d,16'h008d,-16'h003f,16'h00ff,-16'h0222,-16'h0165,16'h00cb,-16'h0076,16'h021b,16'h0004,-16'h00c5,-16'h0097,16'h004d,-16'h003e,-16'h0003,16'h006b,-16'h002e,16'h0039,-16'h0009,16'h00d6,-16'h0028,16'h0048,16'h003b,16'h0055,-16'h006a,-16'h0103,-16'h026d,-16'h00b9,-16'h0062,16'h013c,-16'h0030,16'h00c7,-16'h000a,16'h0048,16'h0127,-16'h0138,-16'h001b,16'h01f7,16'h014b,16'h0006,-16'h003a,-16'h00d1,16'h01ed,16'h0052,16'h003f,-16'h02f3,16'h00ab,16'h005d,16'h0018,16'h00c3,-16'h016d,-16'h00be,16'h000a,16'h00f0,-16'h0084,16'h008f,16'h0171,16'h0091,-16'h00ed,16'h000c,-16'h009c,-16'h0123,16'h00a3,16'h0185,16'h005d,16'h0076,16'h0061,-16'h0031,-16'h013c,-16'h00a0,16'h0139,-16'h00f2,16'h0283,16'h00c3,-16'h013d,-16'h0082,16'h003e,16'h004c,-16'h0011,16'h0086,-16'h0077,16'h007d,16'h0046,16'h00b2,-16'h008a,16'h00db,16'h0000,16'h0036,-16'h012c,-16'h0054,-16'h02fe,-16'h005c,-16'h001a,16'h00bd,-16'h0126,16'h0095,-16'h0019,16'h006a,16'h0164,-16'h02b3,-16'h0027,16'h01f5,16'h0131,-16'h002a,16'h000b,-16'h01f2,16'h01d1,16'h0063,16'h00a7,-16'h0345,16'h004e,16'h0063,-16'h002e,16'h0093,-16'h00ea,-16'h00c8,16'h0032,16'h001b,-16'h0002,16'h0091,16'h0101,16'h0012,-16'h011f,-16'h0042,-16'h010d,-16'h0107,16'h0077,16'h0196,16'h00f1,16'h000e,16'h00bc,-16'h010c,-16'h006f,16'h001c,16'h00de,-16'h008a,16'h0250,-16'h0032,-16'h0153,-16'h00be,16'h000f,16'h002e,16'h001c,16'h007e,-16'h00cf,16'h0083,16'h0095,-16'h0057,-16'h0056,16'h0071,-16'h0028,16'h0036,-16'h00c3,16'h002d,-16'h038d,-16'h0013,-16'h0030,16'h012e,-16'h0086,16'h0142,-16'h009e,-16'h000c,16'h0155,-16'h02b4,-16'h0069,16'h01f7,16'h0199,-16'h0022,-16'h0059,-16'h025d,16'h0228,16'h007c,16'h00d7,-16'h03b0,-16'h0013,16'h00c8,-16'h0004,-16'h0047,-16'h00d5,-16'h0092,16'h001e,16'h0047,-16'h0098,16'h00b0,16'h0163,-16'h014c,-16'h0024,-16'h0061,-16'h008c,-16'h002f,16'h009f,16'h016f,16'h0090,16'h0046,16'h008f,-16'h0142,-16'h0038,-16'h0016,-16'h00d8,-16'h0018,16'h0176,16'h0011,-16'h0104,-16'h012c,16'h007d,16'h0054,-16'h0011,16'h00d5,-16'h002a,16'h007b,16'h005f,16'h002f,-16'h009e,16'h0092,-16'h00e7,16'h008f,-16'h0045,16'h000a,-16'h03d6,16'h0060,16'h0027,16'h00ce,-16'h0063,16'h0178,-16'h0121,-16'h009c,16'h0207,-16'h0280,-16'h001a,16'h022a,16'h011b,-16'h0096,-16'h0026,-16'h0353,16'h0230,16'h0037,16'h006b,-16'h0524,-16'h00b6,16'h00cc,-16'h0020,-16'h006a,-16'h00ae,-16'h003c,-16'h0056,16'h000a,-16'h0056,-16'h0005,16'h016a,-16'h0168,-16'h0004,16'h0006,-16'h0169,16'h004a,16'h006b,16'h01b3,-16'h007e,16'h00d4,16'h006d,-16'h0031,16'h0022,16'h0011,-16'h027c,-16'h010c,16'h0174,16'h0009,-16'h00ee,-16'h013a,-16'h001f,16'h0071,-16'h001a,16'h0088,16'h0019,16'h0072,-16'h0032,-16'h0013,-16'h0124,16'h00dd,-16'h00c1,16'h0029,16'h00a7,16'h009c,-16'h0362,-16'h000b,16'h00e8,16'h0062,-16'h0071,16'h0095,-16'h00f9,-16'h0036,16'h00da,-16'h0269,-16'h0058,16'h0262,16'h009d,-16'h009d,16'h005d,-16'h03f9,16'h028e,-16'h0003,16'h0130,-16'h0551,-16'h0042,16'h0032,16'h0061,16'h00d0,-16'h005c,-16'h0023,-16'h00a3,16'h00af,-16'h005f,16'h0034,16'h018e,-16'h0089,-16'h0050,16'h007b,-16'h0176,16'h00ec,16'h0036,16'h0199,-16'h01ce,16'h00d9,16'h00cd,16'h006a,-16'h00ed,16'h0027,-16'h01da,-16'h0112,16'h0193,-16'h0024,-16'h002e,-16'h0195,-16'h005c,16'h0113,-16'h00a1,16'h0071,-16'h0025,16'h0075,-16'h0054,16'h005e,-16'h0105,16'h004b,-16'h0063,-16'h000b,16'h0064,-16'h003c,-16'h034b,-16'h0020,16'h00ef,16'h0094,-16'h00e2,-16'h0018,-16'h015e,-16'h002b,16'h0078,-16'h0255,16'h001e,16'h028b,16'h00ba,-16'h0066,16'h00b4,-16'h04ef,16'h01f7,-16'h00e0,16'h00f5,-16'h064c,16'h0048,16'h009b,16'h0044,16'h00ee,16'h0017,-16'h0092,16'h0036,16'h0047,16'h001e,-16'h0006,16'h01b8,-16'h00ea,-16'h00a4,16'h001c,-16'h0178,16'h00f8,-16'h0042,16'h00b8,-16'h0241,16'h0047,16'h0057,16'h0002,-16'h00c0,-16'h00c2,-16'h0130,-16'h009f,16'h010a,-16'h0037,-16'h000f,-16'h0269,-16'h00e0,16'h00d7,-16'h0107,16'h0067,-16'h0021,16'h00a5,-16'h009f,16'h007f,-16'h00f4,16'h0067,-16'h006b,-16'h0008,16'h00cc,16'h002e,-16'h0235,16'h0050,16'h00a1,-16'h002a,-16'h0052,16'h002a,-16'h0138,16'h0084,16'h0052,-16'h02a3,-16'h0071,16'h0280,16'h00ad,-16'h0084,16'h0149,-16'h0526,16'h01db,-16'h003d,16'h00e1,-16'h0755,16'h003a,16'h007a,-16'h0010,16'h00a4,16'h009f,-16'h009c,16'h000b,16'h00a9,16'h008b,-16'h0030,16'h013e,-16'h005e,-16'h0142,16'h0026,-16'h0195,16'h0115,-16'h0099,-16'h004a,-16'h01a9,16'h004d,16'h0011,-16'h0066,16'h000c,-16'h0118,-16'h0083,-16'h003c,16'h00b3,-16'h0098,-16'h00bf,-16'h014d,-16'h00ad,16'h0083,-16'h00fc,16'h00a9,-16'h0051,16'h0080,-16'h00e6,16'h00c8,-16'h00f6,-16'h000a,-16'h006d,-16'h00be,16'h0000,-16'h004b,-16'h00c2,16'h006a,16'h00dd,-16'h0020,-16'h00b3,-16'h0078,-16'h00c7,16'h007b,16'h00a5,-16'h0254,-16'h0020,16'h01fc,16'h00a2,-16'h00b2,16'h0095,-16'h04e3,16'h01a5,16'h001f,16'h018a,-16'h07c3,-16'h0068,-16'h001b,-16'h0013,16'h003d,16'h00b7,-16'h0022,16'h00e9,16'h005e,16'h00be,16'h0076,16'h018d,16'h00a1,-16'h0187,16'h0097,-16'h01bb,16'h013a,-16'h0052,-16'h0075,-16'h0109,16'h0034,16'h0086,-16'h009b,16'h006f,-16'h0095,16'h00f0,-16'h0087,16'h0060,-16'h00b0,-16'h007f,-16'h00ae,-16'h004c,16'h00c3,-16'h00ed,16'h010e,-16'h001c,16'h00fe,-16'h00a3,16'h0110,-16'h00c6,-16'h001b,-16'h004a,-16'h001b,-16'h0196,-16'h0024,16'h00a1,16'h0014,16'h00c8,-16'h0025,-16'h011c,-16'h0058,-16'h0067,16'h008c,16'h00c9,-16'h021e,-16'h000e,16'h01ef,16'h0097,-16'h000b,16'h000d,-16'h0584,16'h019f,-16'h0058,16'h00ff,-16'h075c,-16'h00d9,-16'h00e5,-16'h0049,16'h0081,16'h0090,-16'h001c,16'h0095,16'h0054,16'h0012,16'h0023,16'h01bf,16'h00ac,-16'h0094,16'h0148,-16'h02b1,16'h005b,-16'h00c4,-16'h0049,16'h0000,16'h001e,16'h005c,-16'h00e1,16'h00da,-16'h00b5,16'h00f6,16'h0018,16'h00bd,-16'h00af,-16'h012e,16'h00af,-16'h00c7,16'h0123,-16'h0069,16'h00b9,-16'h0062,16'h0139,-16'h0096,16'h0148,-16'h0057,-16'h002e,-16'h004c,-16'h0018,-16'h025a,-16'h00b8,16'h0032,16'h004a,16'h0026,16'h0020,-16'h0130,-16'h001b,16'h000c,16'h001a,16'h00fb,-16'h0218,-16'h0061,16'h0196,16'h00f5,-16'h0051,-16'h0039,-16'h05c4,16'h0129,-16'h0028,16'h00d3,-16'h06c1,-16'h00bd,-16'h007e,-16'h00cc,-16'h0034,16'h0117,16'h004a,16'h0071,16'h00ab,-16'h006d,16'h0037,16'h0159,16'h006d,16'h000c,16'h0179,-16'h0281,-16'h017e,-16'h00c6,-16'h0022,16'h001a,16'h00d3,16'h0024,-16'h0165,16'h0070,-16'h00f3,16'h00fb,16'h0028,16'h0103,-16'h0093,-16'h0073,16'h0171,-16'h0032,16'h0119,-16'h011e,16'h00f9,16'h0017,16'h0109,-16'h005c,16'h00b5,-16'h0061,16'h002f,-16'h011f,16'h007b,-16'h021c,-16'h0146,-16'h0035,16'h0089,16'h008d,16'h0020,-16'h00aa,16'h002e,16'h0009,-16'h0092,16'h015e,-16'h01f3,-16'h0068,16'h0103,16'h010b,-16'h008f,-16'h001c,-16'h0644,16'h00b1,-16'h0048,16'h0078,-16'h0610,-16'h0039,-16'h003a,-16'h009c,16'h001b,16'h00cc,16'h0049,16'h0040,16'h0089,-16'h003d,16'h0043,16'h014a,16'h00fb,-16'h007d,16'h0188,-16'h020f,-16'h0030,16'h0039,-16'h00c7,16'h0091,16'h0083,-16'h004f,-16'h0089,16'h0044,-16'h010d,-16'h0005,16'h0082,16'h013b,-16'h0053,16'h0092,16'h01cc,-16'h0053,16'h001a,-16'h0276,16'h0065,-16'h0092,16'h0107,-16'h006f,16'h00cc,-16'h0019,16'h003a,-16'h00fc,-16'h0046,-16'h006c,-16'h019e,16'h0075,-16'h0011,-16'h0020,16'h009f,-16'h006d,-16'h0055,-16'h000d,-16'h0072,16'h012b,-16'h00f6,-16'h00bf,16'h01a6,16'h00e9,-16'h007b,16'h0063,-16'h06b6,16'h0028,-16'h00a6,16'h0090,-16'h052f,16'h0005,16'h0001,-16'h0073,16'h0060,16'h015d,16'h00b0,-16'h002f,16'h0092,16'h000b,-16'h005c,16'h017a,16'h00a1,16'h0007,16'h0108,-16'h02a9,-16'h001c,16'h00c8,-16'h01d3,16'h0067,16'h009b,-16'h0039,16'h0001,-16'h0094,-16'h0078,-16'h00bf,-16'h0003,16'h0096,-16'h003e,16'h0150,16'h017b,-16'h003b,16'h0008,-16'h042a,16'h00ce,-16'h00a1,16'h005d,-16'h00bd,16'h009a,16'h000b,-16'h0028,-16'h00e8,-16'h00c0,16'h009f,-16'h00fd,16'h00c3,16'h00d5,16'h0083,-16'h0046,-16'h00da,16'h0061,16'h0056,16'h004f,16'h0153,-16'h0031,-16'h016c,16'h0162,16'h0123,-16'h0027,16'h00b1,-16'h0652,16'h0098,-16'h0114,16'h008e,-16'h048e,16'h0012,16'h005d,-16'h0027,16'h009f,16'h0123,16'h007d,-16'h00ac,16'h00ef,-16'h0003,-16'h0122,16'h00d8,16'h006d,16'h00e6,16'h00d7,-16'h0330,16'h0063,16'h00f7,-16'h029f,16'h0084,16'h0064,16'h0027,16'h0079,-16'h006b,-16'h000c,-16'h01f8,-16'h0059,16'h00d9,-16'h0046,16'h010f,16'h014b,-16'h0050,16'h001b,-16'h04ab,16'h0089,-16'h00bb,-16'h0043,-16'h0108,16'h00c2,16'h0047,16'h0058,-16'h004a,-16'h0084,16'h0116,-16'h00dc,16'h011b,16'h012a,-16'h00b5,-16'h0009,-16'h0047,16'h0050,16'h0069,16'h004d,16'h0184,-16'h0070,-16'h019c,16'h016d,16'h0123,-16'h0010,16'h00b4,-16'h0538,16'h0086,-16'h0163,16'h0064,-16'h0422,16'h0030,16'h011d,-16'h0066,16'h0103,16'h0150,16'h0064,-16'h005f,16'h0148,-16'h0047,-16'h0141,16'h00cb,16'h0004,16'h00a0,-16'h02e2,-16'h02da,16'h0005,16'h019c,-16'h0330,-16'h002a,16'h0090,16'h008a,16'h01dc,-16'h006c,16'h00d7,-16'h0195,-16'h008a,16'h0023,16'h004f,16'h0114,16'h012b,-16'h0094,16'h0010,-16'h0528,16'h006d,-16'h0056,-16'h0041,-16'h014d,16'h00b9,16'h00e9,-16'h0053,16'h005d,-16'h0050,16'h00de,-16'h0004,16'h017c,16'h00ae,-16'h01a5,16'h0041,16'h001e,-16'h005b,16'h00fa,-16'h005e,16'h0102,-16'h0019,-16'h01da,16'h0146,16'h006e,-16'h0081,16'h00b1,-16'h03ca,16'h0127,-16'h008c,16'h0016,-16'h03d9,16'h0093,16'h003c,16'h0018,16'h00bd,16'h012f,16'h0015,16'h006b,16'h0104,-16'h008d,-16'h022a,16'h007b,-16'h0086,-16'h0039,-16'h07ea,-16'h030d,16'h0037,16'h0132,-16'h0299,-16'h0112,16'h0009,16'h00e8,16'h01e5,-16'h003b,16'h0108,-16'h00a0,-16'h0036,16'h0021,16'h000d,16'h00a8,16'h0116,-16'h017e,-16'h0036,-16'h0370,16'h000f,-16'h0104,16'h0063,-16'h0132,16'h00f0,16'h017d,-16'h0043,16'h0089,16'h0005,16'h0018,16'h0079,16'h01d8,16'h0019,-16'h042f,16'h00a8,-16'h0024,-16'h0057,16'h008c,-16'h01a1,16'h0184,16'h0034,-16'h01dd,16'h0120,16'h007a,-16'h00c8,16'h0062,-16'h02a9,16'h00d1,-16'h0047,16'h007a,-16'h039d,16'h002e,16'h00e9,-16'h0038,16'h0024,16'h01e3,16'h0023,16'h000e,-16'h002e,-16'h008b,-16'h033a,16'h0170,-16'h00af,-16'h00b0,-16'h0881,-16'h02d8,16'h00ac,16'h00e6,-16'h01ef,-16'h0155,16'h004d,16'h01ae,16'h01ed,-16'h002a,16'h011e,16'h00a1,-16'h0055,16'h00aa,16'h00aa,16'h0160,16'h00d2,-16'h0073,-16'h001a,-16'h025d,-16'h001b,-16'h0158,16'h0004,-16'h00b5,16'h01bd,16'h0131,16'h0005,-16'h005a,16'h0002,-16'h00d4,16'h0094,16'h01b2,16'h00b8,-16'h069f,16'h0083,16'h0020,-16'h0025,16'h0121,-16'h0273,16'h00fa,16'h00d3,-16'h013b,16'h012e,-16'h0013,-16'h006d,-16'h003b,-16'h0242,16'h010d,16'h0022,16'h0068,-16'h0311,16'h009a,16'h0092,-16'h00ff,-16'h00f7,16'h015c,-16'h0047,-16'h009e,-16'h00cb,-16'h001c,-16'h0343,16'h01a4,-16'h009b,-16'h011c,-16'h04bc,-16'h02b6,16'h00bd,16'h0003,-16'h015d,-16'h0197,16'h0109,16'h0152,16'h0268,16'h0032,16'h010a,16'h00f9,-16'h003e,16'h00c4,16'h00ab,16'h00ae,16'h00d7,-16'h004b,16'h002b,-16'h01be,16'h0006,-16'h0199,-16'h0053,16'h0068,16'h015e,16'h00f6,-16'h0087,16'h0019,-16'h0030,-16'h0117,16'h00ab,16'h018e,-16'h0013,-16'h04db,16'h00d9,16'h000f,-16'h006e,-16'h0022,-16'h021c,16'h0166,16'h0070,-16'h0065,16'h012f,16'h0006,-16'h0057,-16'h00b0,-16'h01ab,16'h006b,16'h0165,16'h008c,-16'h0328,16'h004a,16'h00d4,-16'h0048,-16'h0052,16'h0189,16'h0012,-16'h0007,-16'h0099,-16'h0059,-16'h032f,16'h0186,16'h0010,-16'h0168,-16'h026f,-16'h01da,16'h00b3,-16'h02b9,-16'h00d8,-16'h0179,16'h00a0,-16'h0022,16'h01c0,16'h0074,16'h00a8,16'h0175,-16'h005c,16'h0107,-16'h0038,16'h0062,16'h0056,16'h006b,16'h0007,-16'h01d3,16'h000f,-16'h0175,-16'h0139,16'h0201,16'h0164,16'h00ed,16'h0034,16'h0043,16'h000f,-16'h0171,-16'h0028,16'h01fe,-16'h0057,-16'h0251,16'h00f7,-16'h0036,-16'h0127,-16'h0015,-16'h0121,16'h0186,16'h00f7,-16'h0073,16'h00ed,-16'h0029,-16'h004b,-16'h0163,-16'h01f0,16'h0011,16'h0261,16'h0014,-16'h02d2,16'h0063,16'h009b,-16'h0148,16'h00b3,16'h017b,-16'h0029,16'h004c,-16'h0163,16'h000c,-16'h0298,16'h014b,-16'h005a,-16'h0144,-16'h0127,-16'h0185,16'h0131,-16'h04c3,-16'h0090,-16'h0195,16'h004a,-16'h0057,16'h01cd,16'h004f,16'h0004,16'h0118,-16'h004d,16'h00d3,-16'h006f,16'h014e,16'h00cb,16'h0089,16'h0044,-16'h0180,16'h0001,-16'h00dd,-16'h00db,16'h0231,16'h0198,16'h00c6,16'h0059,16'h00cd,-16'h0011,-16'h00fd,-16'h0096,16'h013e,-16'h0055,-16'h0161,16'h000d,-16'h004e,-16'h00c8,-16'h004c,-16'h00ae,16'h0165,16'h0038,-16'h004b,-16'h0014,-16'h002d,16'h0018,-16'h01a1,-16'h0159,-16'h00c6,16'h026c,16'h0051,-16'h021c,16'h00ea,16'h0029,-16'h010f,16'h00e7,16'h01dc,16'h0030,16'h007d,-16'h016d,-16'h0036,-16'h0166,16'h013f,-16'h0007,-16'h0133,-16'h000e,-16'h0091,16'h0182,-16'h03d8,16'h0004,-16'h01f5,16'h0090,-16'h00db,16'h005e,16'h005f,-16'h0025,16'h00d7,-16'h0078,16'h00b6,-16'h002f,16'h01b4,-16'h001b,16'h008b,16'h009c,-16'h00e3,16'h0056,-16'h004e,-16'h0081,16'h01ab,16'h013c,16'h001b,-16'h0050,16'h00ca,16'h00a9,-16'h0037,-16'h007b,16'h0126,-16'h0043,16'h0002,-16'h008a,16'h000d,16'h0022,-16'h009f,-16'h009b,16'h012b,16'h0008,-16'h017d,-16'h0035,-16'h0024,16'h00fe,-16'h010f,-16'h0199,-16'h00c0,16'h0276,16'h00db,-16'h00c7,-16'h0045,16'h0060,-16'h0104,16'h0158,16'h023d,16'h002b,16'h008a,-16'h00a8,16'h006e,-16'h00d0,16'h0149,-16'h003e,-16'h00a6,16'h004e,16'h000b,16'h012f,-16'h026e,-16'h003d,-16'h01a7,16'h0056,-16'h0029,-16'h00d7,16'h001e,-16'h0049,16'h0121,-16'h0005,16'h0106,-16'h0039,16'h02a8,-16'h005e,16'h0067,16'h0038,-16'h0118,16'h002e,-16'h0029,-16'h004b,16'h00f7,16'h0183,-16'h007f,-16'h0125,16'h00e6,16'h00ac,-16'h00e8,-16'h00d5,16'h0127,16'h0092,-16'h0022,-16'h011e,-16'h00bb,16'h0102,16'h010f,16'h003b,16'h00c4,16'h0033,-16'h0113,16'h010d,16'h00ea,-16'h0069,16'h0162,16'h0138,16'h004e,16'h017c,-16'h00f2,16'h0039,-16'h0091,-16'h0051,16'h0136,-16'h0046,-16'h0057,-16'h00b7,-16'h00ca,-16'h00d6,16'h00a4,16'h0112,-16'h00b0,-16'h000c,-16'h0150,16'h007c,-16'h0021,16'h00e0,-16'h009d,16'h01d6,16'h00d0,-16'h0038,16'h0054,16'h0004,-16'h0055,16'h0171,-16'h005d,16'h0019,16'h01b8,-16'h0056,-16'h0012,16'h003e,-16'h0020,16'h0008,16'h00ad,-16'h002d,16'h007f,16'h014c,-16'h005a,16'h0198,16'h0043,16'h0063,16'h009f,-16'h00fb,-16'h009b,-16'h014f,-16'h0044,-16'h00c8,-16'h0099,16'h00b8,-16'h005f,16'h00c8,16'h00b6,-16'h0004,16'h0094,-16'h0027,-16'h0170,16'h0144,16'h00ab,-16'h0082,16'h0111,16'h0130,16'h006d,16'h01da,-16'h00c7,16'h0053,16'h0015,16'h0063,16'h00f9,16'h0060,16'h0032,-16'h007b,-16'h0138,-16'h016e,16'h00b7,16'h00da,-16'h0070,-16'h0005,-16'h0174,16'h003f,16'h0019,16'h009c,-16'h0074,16'h01f6,16'h018d,16'h0015,-16'h000d,16'h0068,-16'h0021,16'h00de,-16'h0077,16'h0037,16'h018b,-16'h0016,-16'h0026,-16'h0014,-16'h0036,-16'h000f,16'h002d,16'h0008,16'h00e0,16'h00b3,-16'h00ec,16'h0104,-16'h002e,16'h0040,16'h013a,-16'h009d,-16'h0041,-16'h0174,-16'h009f,-16'h0141,-16'h0001,16'h00c5,16'h003d,16'h00a2,16'h0111,16'h002f,16'h0082,16'h002c,-16'h0136,16'h01f7,16'h0074,-16'h0096,16'h0109,16'h00ff,16'h0061,16'h0275,-16'h0198,16'h00d9,-16'h0021,16'h0042,16'h0085,16'h0018,-16'h006c,-16'h0074,-16'h0143,-16'h00de,16'h006b,16'h00ad,-16'h003d,16'h004a,-16'h0235,16'h006a,-16'h005e,16'h009d,16'h0079,16'h02a4,16'h01bc,16'h007a,-16'h0083,16'h0030,-16'h005c,16'h00ec,-16'h0095,-16'h008d,16'h0184,-16'h0084,-16'h0005,-16'h00e9,16'h0030,16'h0025,16'h008a,16'h0001,16'h009c,16'h00b7,-16'h00c2,16'h0093,-16'h0031,-16'h001f,16'h01be,16'h000a,16'h0069,-16'h00c1,-16'h00a6,-16'h008f,16'h0012,16'h0095,16'h001d,16'h0042,16'h014e,16'h0030,16'h006f,-16'h0044,-16'h012b,16'h01b4,16'h001f,-16'h0070,16'h00ae,16'h000d,16'h0089,16'h022e,-16'h018c,-16'h0028,16'h0019,-16'h0002,-16'h0002,16'h0010,-16'h0082,-16'h007b,-16'h0138,-16'h0082,-16'h002a,16'h0023,16'h0005,-16'h001b,-16'h0191,16'h003c,-16'h0040,16'h0080,16'h0036,16'h032f,16'h0208,-16'h001b,-16'h00af,16'h009e,-16'h0067,16'h00b2,-16'h0034,-16'h0088,16'h0184,-16'h0148,-16'h004d,-16'h0121,16'h000b,-16'h010a,16'h0058,16'h000a,16'h004f,16'h009d,-16'h0158,16'h0094,-16'h0052,-16'h0034,16'h012b,16'h0034,16'h00a8,-16'h0109,-16'h011c,-16'h00bd,16'h0034,16'h0049,-16'h0041,16'h00be,16'h00ee,16'h003c,16'h00bc,-16'h007c,-16'h0090,16'h01ac,16'h007e,-16'h0024,16'h00ea,-16'h0099,16'h00c6,16'h0231,-16'h0123,-16'h01cf,-16'h000f,-16'h0035,16'h0015,16'h0048,-16'h0170,-16'h0053,-16'h0127,16'h0059,-16'h011d,16'h0041,16'h0079,16'h0038,-16'h017e,16'h0000,16'h0000,-16'h0014,16'h0076,16'h01e9,16'h00f3,16'h003a,-16'h0182,16'h0146,-16'h0088,-16'h0047,-16'h0063,-16'h00d9,16'h01fd,-16'h0179,-16'h009a,-16'h012e,16'h003e,-16'h00e7,16'h0083,-16'h0003,-16'h009b,16'h0070,-16'h0163,16'h0093,-16'h0049,16'h0019,16'h00be,16'h0003,16'h0044,-16'h011e,-16'h01c0,-16'h0037,16'h0008,16'h009e,-16'h0015,16'h00e7,16'h0066,16'h00a3,16'h015a,-16'h006f,16'h006b,16'h019d,16'h007c,16'h0037,16'h0049,-16'h0146,16'h00c7,16'h01ee,-16'h00ae,-16'h0317,16'h006c,16'h0013,16'h000a,16'h0092,-16'h01fa,16'h004a,-16'h0077,16'h00ed,-16'h015d,-16'h0009,16'h0055,16'h0129,-16'h005b,-16'h000d,16'h0000,-16'h007b,16'h00f5,16'h0226,16'h00ea,16'h002a,-16'h00d0,16'h01b5,-16'h0123,-16'h00fe,16'h0029,-16'h0090,16'h020f,-16'h0151,-16'h00a3,-16'h00ea,16'h0064,-16'h00dd,16'h0064,16'h005f,-16'h00f6,16'h003f,-16'h00d5,16'h00ba,-16'h0087,-16'h0045,16'h0079,16'h0019,16'h008c,-16'h00e4,-16'h0268,16'h0016,-16'h0044,16'h00cf,16'h0052,16'h00ba,16'h009c,16'h0030,16'h00fd,-16'h019a,16'h00c0,16'h018e,16'h0072,-16'h0030,-16'h000e,-16'h01ba,16'h00cc,16'h012c,-16'h00c2,-16'h0350,16'h0054,16'h003e,16'h0010,16'h0015,-16'h01de,-16'h002f,16'h0017,16'h0167,-16'h00a9,16'h00b3,16'h00bc,16'h011e,-16'h00f4,-16'h0043,-16'h002f,-16'h00bc,16'h0112,16'h011f,-16'h0050,16'h0011,-16'h008f,16'h01a1,-16'h01df,-16'h00c4,16'h00d3,-16'h0116,16'h0244,16'h0060,-16'h0080,-16'h0117,16'h0054,-16'h0088,16'h0008,16'h0077,-16'h0100,16'h0016,16'h005c,16'h011e,16'h0000,-16'h0036,-16'h002d,16'h0061,16'h00b9,-16'h011b,-16'h03c3,-16'h0054,16'h0013,16'h0146,-16'h001d,16'h00a9,16'h0007,16'h0010,16'h019a,-16'h02a6,16'h00d6,16'h01f3,16'h0138,16'h0050,-16'h0030,-16'h02a5,16'h0136,16'h00c6,-16'h000a,-16'h0479,16'h0031,16'h00d5,-16'h004e,-16'h0025,-16'h01c7,-16'h005c,-16'h00a7,16'h0147,-16'h00bb,16'h0059,16'h0112,16'h0088,-16'h00bc,-16'h0025,-16'h002e,-16'h0187,16'h010a,16'h015d,-16'h0066,16'h00a7,-16'h000a,16'h0107,-16'h0143,-16'h0107,16'h00cc,-16'h012d,16'h01ed,16'h006b,-16'h012e,-16'h00e0,-16'h0030,16'h0054,-16'h0014,-16'h0017,-16'h00df,16'h009c,16'h0058,16'h00df,-16'h000c,16'h0024,-16'h00da,16'h0010,16'h0006,-16'h010b,-16'h045f,-16'h001e,16'h0003,16'h012f,-16'h0078,16'h0120,-16'h0029,16'h0036,16'h0137,-16'h03b2,16'h005f,16'h011d,16'h014e,16'h000b,-16'h0087,-16'h038b,16'h016e,16'h00de,16'h0080,-16'h0628,16'h006c,16'h0084,-16'h0004,-16'h0026,-16'h01fd,-16'h0084,-16'h000e,16'h00c9,-16'h0002,16'h00c9,16'h00e3,-16'h000b,-16'h0059,-16'h004d,-16'h00a1,-16'h0116,16'h0055,16'h0101,-16'h0010,-16'h0016,16'h0017,-16'h007a,-16'h0050,-16'h000f,-16'h000b,-16'h0077,16'h022c,16'h00d9,-16'h0149,-16'h0080,-16'h0022,16'h004e,16'h009a,16'h003f,-16'h0081,16'h0045,16'h007e,16'h005b,-16'h0048,16'h0060,-16'h00ea,-16'h0064,16'h0054,-16'h0079,-16'h042b,16'h00c1,16'h00fa,16'h00d5,-16'h00d3,16'h00b3,-16'h0062,16'h002b,16'h0159,-16'h0485,16'h0099,16'h0149,16'h020f,-16'h001e,-16'h0084,-16'h0405,16'h01ae,16'h007c,16'h0096,-16'h082c,16'h008b,16'h00c1,16'h006b,-16'h016e,-16'h01c1,-16'h0081,16'h0073,-16'h0001,16'h000f,16'h00d3,16'h00ed,-16'h01d9,16'h0017,-16'h0011,-16'h0070,-16'h00b3,16'h004f,16'h00ea,16'h002f,16'h002d,16'h006c,-16'h00d0,16'h00d4,16'h0002,-16'h00d7,-16'h007a,16'h0194,16'h006a,-16'h004f,-16'h00f5,-16'h001a,16'h0076,16'h0044,16'h00aa,-16'h002f,-16'h0016,16'h00cb,16'h00b3,-16'h0030,16'h005a,-16'h010e,-16'h002a,16'h0038,-16'h0057,-16'h03bb,16'h0074,16'h0080,16'h009d,-16'h00e1,16'h00b4,-16'h00d4,-16'h005c,16'h015f,-16'h040c,16'h00ed,16'h00e3,16'h0133,-16'h0009,-16'h00a9,-16'h0379,16'h019c,16'h00a3,16'h007d,-16'h08ea,-16'h0056,16'h00cf,16'h0053,-16'h0092,-16'h01fe,16'h004d,-16'h00ef,16'h0079,16'h001a,16'h0054,16'h00e0,-16'h016e,16'h00ba,16'h0050,-16'h00ae,16'h0069,-16'h0025,16'h0009,-16'h0083,16'h00ce,16'h00a8,-16'h0039,16'h0025,-16'h0013,-16'h01b8,-16'h0061,16'h0167,-16'h0015,-16'h009d,-16'h0165,16'h003f,-16'h0003,16'h0040,16'h00b9,16'h002e,-16'h0024,16'h00a7,16'h007a,-16'h0097,16'h00cf,-16'h0074,16'h0000,16'h00d9,-16'h00c5,-16'h03f6,16'h00b0,16'h00e8,16'h0093,-16'h00b0,16'h00cf,-16'h0067,-16'h00f0,16'h0131,-16'h03e0,16'h0102,16'h012a,16'h011b,-16'h0040,16'h005b,-16'h03f2,16'h01d7,-16'h0065,16'h00c8,-16'h0a01,-16'h003c,16'h0065,16'h008b,16'h008f,-16'h0187,16'h0058,-16'h00ba,16'h0091,-16'h0006,-16'h0031,16'h011c,-16'h009d,16'h00c0,16'h0043,-16'h0106,16'h009b,-16'h0083,16'h0033,-16'h0169,16'h00b8,16'h008c,16'h001e,-16'h00da,-16'h000f,-16'h0122,-16'h0048,16'h0188,16'h0071,16'h0050,-16'h0132,-16'h000b,16'h008d,16'h001a,16'h00c7,-16'h0057,-16'h0024,-16'h00e0,16'h006b,-16'h00b2,16'h00dd,-16'h0051,-16'h0076,16'h00c0,-16'h00a1,-16'h03f7,16'h0045,16'h008b,16'h0019,-16'h00be,-16'h0078,-16'h0026,-16'h009f,16'h00bf,-16'h039f,16'h00c9,16'h0125,16'h00c5,-16'h007c,16'h015c,-16'h031d,16'h01a9,-16'h00bb,16'h011f,-16'h098f,-16'h0005,16'h0012,16'h0076,16'h011b,-16'h0148,16'h005f,16'h0072,16'h006c,16'h000b,16'h0006,16'h008c,-16'h0084,-16'h0015,16'h000d,-16'h0176,16'h0138,-16'h00a6,-16'h0014,-16'h01ab,16'h00c6,-16'h0044,-16'h0016,-16'h00f4,-16'h00a6,-16'h0101,-16'h004e,16'h01ee,16'h000b,16'h0049,-16'h0194,-16'h0096,16'h00a5,16'h002a,16'h0060,-16'h006f,16'h0049,-16'h00b3,16'h009a,-16'h00a5,16'h008c,-16'h00c1,-16'h0057,16'h0054,-16'h0100,-16'h0484,16'h004d,16'h00fb,-16'h0005,-16'h0059,-16'h00b1,-16'h0082,-16'h003a,16'h00f3,-16'h0356,-16'h000d,16'h01bd,16'h00d2,-16'h006a,16'h010b,-16'h027b,16'h0135,-16'h0030,16'h0112,-16'h0856,-16'h002a,16'h0023,16'h005e,16'h00ba,-16'h00ea,16'h0029,16'h0101,16'h005c,16'h00a9,16'h0007,16'h00fa,16'h000c,-16'h0104,16'h000b,-16'h0122,16'h00fa,-16'h0099,-16'h009c,-16'h00d3,16'h0095,-16'h000a,-16'h002b,16'h0000,-16'h0161,-16'h00ae,16'h0033,16'h0160,-16'h0055,-16'h0015,-16'h013f,-16'h0071,16'h006b,-16'h010f,16'h0047,-16'h004c,16'h009e,-16'h0058,16'h0117,-16'h0093,16'h00b4,-16'h00a7,-16'h002a,-16'h0005,-16'h008e,-16'h0337,-16'h0039,16'h0051,-16'h003c,-16'h0058,-16'h003d,16'h0014,16'h0087,16'h00e9,-16'h02dc,16'h0000,16'h0182,16'h010e,-16'h00b5,16'h00e0,-16'h0244,16'h0158,16'h002c,16'h00f2,-16'h084b,-16'h00a8,-16'h0067,-16'h001e,16'h0071,-16'h007f,16'h0014,16'h0068,16'h0073,16'h00a8,-16'h0089,16'h0128,16'h00bf,-16'h00b0,16'h007f,-16'h0149,16'h0128,-16'h00b3,-16'h0102,-16'h0010,16'h008c,16'h0036,-16'h0054,16'h00b2,-16'h00bc,16'h0103,16'h0000,16'h0125,-16'h006d,-16'h0086,-16'h0015,-16'h0037,16'h007e,-16'h0083,16'h005e,-16'h00a7,16'h0118,-16'h0155,16'h016a,-16'h000d,16'h000c,-16'h007f,-16'h0050,-16'h0143,-16'h004b,-16'h01b5,-16'h004b,16'h0060,-16'h003f,-16'h0098,-16'h001f,-16'h000e,16'h004e,16'h016d,-16'h0176,-16'h0028,16'h0177,16'h0141,16'h004a,16'h0052,-16'h02ee,16'h018c,16'h003b,16'h0091,-16'h0849,-16'h00e6,-16'h0013,-16'h0004,16'h0005,-16'h0075,16'h0023,16'h007a,16'h003e,16'h005a,16'h0037,16'h0117,16'h0128,-16'h006a,16'h00d5,-16'h01ef,16'h002b,-16'h009d,-16'h00b0,16'h0067,16'h00a2,-16'h002a,-16'h0141,16'h0098,-16'h00dd,16'h0134,16'h004b,16'h018f,-16'h0046,-16'h0070,16'h0172,-16'h0067,16'h00ef,-16'h011c,16'h00ba,-16'h00cf,16'h0111,-16'h0104,16'h010f,16'h0035,16'h001e,-16'h005a,16'h0097,-16'h0212,-16'h0071,-16'h0171,16'h0031,-16'h0010,-16'h0085,-16'h00fe,16'h000b,16'h006c,16'h002f,16'h015f,-16'h011f,-16'h0033,16'h0152,16'h00f9,16'h001d,16'h0042,-16'h03bb,16'h009b,-16'h0025,16'h0079,-16'h08b8,-16'h0092,-16'h0070,-16'h0050,-16'h001c,-16'h0091,-16'h0033,-16'h004e,16'h0072,16'h004f,-16'h0009,16'h0132,16'h0124,-16'h0073,16'h0119,-16'h01cd,-16'h019c,-16'h009d,-16'h00a4,16'h0041,16'h00d8,-16'h006b,-16'h007c,16'h0128,-16'h0155,16'h0168,16'h006f,16'h01a8,-16'h0061,-16'h001d,16'h0190,-16'h0016,16'h00b6,-16'h020c,16'h006f,-16'h0075,16'h014c,-16'h009d,16'h00f4,16'h00bb,16'h0041,-16'h00d9,16'h0015,-16'h011d,-16'h00b1,-16'h0159,-16'h001f,-16'h004c,16'h0027,-16'h0056,16'h0029,16'h0015,16'h006e,16'h018c,-16'h01d0,-16'h00f1,16'h017d,16'h0112,16'h0096,16'h0038,-16'h045a,-16'h0059,16'h0030,16'h001a,-16'h084d,-16'h0008,-16'h004b,16'h0012,16'h0015,-16'h0050,-16'h000c,-16'h00b9,16'h0078,-16'h000b,-16'h0046,16'h0130,16'h0121,-16'h0064,16'h00c6,-16'h0119,-16'h00b3,16'h0056,-16'h0115,16'h0031,16'h00e2,-16'h00ea,16'h0039,16'h00aa,-16'h008f,16'h005c,16'h00fd,16'h01b8,-16'h0058,16'h00f6,16'h0161,16'h0021,16'h00e6,-16'h030d,16'h0075,-16'h0071,16'h00a3,-16'h00de,16'h0157,16'h0088,-16'h0014,-16'h0174,-16'h000c,16'h0013,-16'h00f5,-16'h0102,16'h000e,-16'h00c1,16'h0044,16'h0000,16'h008c,-16'h0028,16'h000c,16'h01b3,-16'h00b6,-16'h005a,16'h0130,16'h0121,-16'h0007,16'h0025,-16'h048e,-16'h0091,-16'h00f5,16'h0059,-16'h07c2,-16'h0065,-16'h0053,-16'h005a,16'h002c,16'h0020,-16'h0034,-16'h0012,16'h00b6,-16'h0028,-16'h00c7,16'h00eb,16'h00e4,16'h0065,16'h00e8,-16'h01b0,-16'h0046,16'h008c,-16'h0248,16'h009f,16'h00fd,-16'h006f,16'h0069,16'h004e,-16'h007c,-16'h0100,16'h005d,16'h019b,-16'h0045,16'h0192,16'h0104,-16'h0011,16'h00c2,-16'h0470,16'h008d,-16'h00fa,16'h0021,-16'h014a,16'h0145,16'h0062,16'h0016,-16'h0170,-16'h0056,16'h0125,-16'h009f,-16'h00c0,16'h0087,-16'h0091,-16'h004c,16'h002c,16'h002f,16'h008e,-16'h0031,16'h0184,-16'h00c5,-16'h00c8,16'h0139,16'h0164,16'h0002,16'h005f,-16'h0408,16'h0000,-16'h0102,16'h00cf,-16'h06de,16'h0058,16'h000c,-16'h009f,16'h0114,16'h0017,-16'h001c,-16'h0090,16'h00f7,16'h003e,-16'h015f,16'h013c,16'h0073,16'h0064,16'h0006,-16'h01b2,-16'h0027,16'h0100,-16'h02bf,16'h001d,16'h00f4,16'h0009,16'h0155,-16'h0032,16'h0019,-16'h0221,16'h0020,16'h017d,-16'h0016,16'h0199,16'h00ef,-16'h000b,16'h0037,-16'h042e,16'h007e,-16'h003e,-16'h0056,-16'h00c8,16'h0130,16'h00b4,-16'h0007,-16'h0160,-16'h00a1,16'h0135,-16'h006d,-16'h0027,16'h00b7,-16'h013c,16'h000e,-16'h0028,16'h0025,16'h00a9,-16'h000a,16'h0144,-16'h0095,-16'h00e6,16'h0133,16'h013f,-16'h002e,16'h007c,-16'h02f7,16'h0054,-16'h009b,16'h008c,-16'h05aa,-16'h003f,16'h0027,-16'h0047,16'h0118,16'h0051,-16'h0065,-16'h005e,16'h01dc,-16'h00a3,-16'h0202,16'h0101,-16'h0031,16'h00eb,-16'h02f9,-16'h02af,16'h0075,16'h00fd,-16'h0260,-16'h00d7,16'h008b,16'h00b2,16'h018a,-16'h0093,16'h008a,-16'h0139,16'h0039,16'h00cf,16'h008b,16'h0161,16'h00fa,-16'h0003,16'h002f,-16'h0322,16'h0082,-16'h0083,-16'h0078,-16'h018b,16'h0152,16'h00af,16'h000b,-16'h00b0,-16'h0093,16'h006c,-16'h000c,16'h006d,16'h0002,-16'h020d,16'h006e,16'h0065,-16'h0004,16'h00ec,-16'h01b1,16'h0179,-16'h004b,-16'h00cc,16'h0186,16'h00c4,-16'h0041,16'h00af,-16'h023e,16'h00ce,-16'h0044,16'h00c5,-16'h04fb,16'h0086,16'h0022,-16'h006a,16'h005e,16'h00a4,-16'h00e8,-16'h006c,16'h01c9,-16'h00b0,-16'h01e4,16'h012f,-16'h0065,16'h0088,-16'h06aa,-16'h0212,16'h0076,16'h00c8,-16'h01c1,-16'h0157,16'h007f,16'h019b,16'h01f3,-16'h0025,16'h00c2,-16'h0014,16'h0001,16'h017e,16'h00e5,16'h0172,16'h00ac,-16'h006d,16'h0049,-16'h02a0,-16'h000c,-16'h00ac,-16'h0027,-16'h012d,16'h012f,16'h011c,-16'h00ab,-16'h0072,-16'h0070,16'h002b,16'h005a,16'h0130,16'h0027,-16'h03cd,16'h0066,16'h006c,-16'h0076,16'h012e,-16'h0228,16'h014e,16'h0107,-16'h006f,16'h016d,16'h0115,-16'h003e,-16'h0001,-16'h01d5,16'h00a0,-16'h005f,16'h0047,-16'h0432,16'h0070,16'h004d,-16'h0103,-16'h0035,16'h00df,-16'h00fe,-16'h0068,16'h00dd,-16'h00b5,-16'h0320,16'h0146,-16'h00cb,-16'h00a5,-16'h06c4,-16'h0271,16'h0097,16'h007b,-16'h00d7,-16'h015b,16'h0055,16'h0201,16'h023a,-16'h0026,16'h00d5,16'h00f4,16'h004a,16'h01a4,16'h00c7,16'h00dd,16'h0037,-16'h0081,16'h002a,-16'h0172,-16'h0079,-16'h00de,16'h0005,-16'h00b3,16'h0165,16'h00d3,-16'h004d,-16'h011b,16'h003c,-16'h00b0,16'h011a,16'h011e,16'h003d,-16'h0591,16'h0093,16'h009a,-16'h0059,16'h00b1,-16'h01b4,16'h0154,16'h0163,-16'h0069,16'h0068,16'h004f,-16'h0059,-16'h00ee,-16'h01c0,16'h0066,16'h0085,16'h0028,-16'h0438,16'h008d,16'h00d9,-16'h011f,-16'h00fa,16'h0140,-16'h004c,-16'h0093,16'h0041,-16'h0057,-16'h0300,16'h01a6,-16'h0013,-16'h013e,-16'h03fd,-16'h02d5,16'h00ae,-16'h002c,-16'h0116,-16'h01a6,16'h009f,16'h016d,16'h01e9,16'h0072,16'h0078,16'h00c1,16'h001e,16'h014a,16'h0047,16'h00af,-16'h005c,16'h0006,16'h0061,-16'h0167,16'h0040,-16'h012a,-16'h00e9,16'h00fe,16'h017b,16'h00ce,-16'h009f,-16'h0106,-16'h003a,-16'h0198,16'h005f,16'h0146,-16'h0033,-16'h03d5,16'h0091,16'h005a,-16'h0084,-16'h0090,-16'h0164,16'h0134,16'h01a2,16'h0025,16'h0111,-16'h005e,16'h000b,-16'h0176,-16'h0198,16'h009f,16'h01b5,16'h007d,-16'h03a9,16'h00a1,16'h001e,-16'h0085,16'h000d,16'h00fc,-16'h004b,-16'h001c,16'h0050,-16'h0083,-16'h028c,16'h0223,16'h0000,-16'h0277,-16'h022a,-16'h0255,16'h0099,-16'h020f,-16'h00ba,-16'h019e,16'h0139,16'h0085,16'h01c7,16'h00e7,16'h0011,16'h010b,16'h002a,16'h0163,-16'h00bd,16'h00f9,16'h0015,16'h00ca,16'h008b,-16'h01bd,16'h002c,-16'h00a3,-16'h00eb,16'h0197,16'h017a,16'h00ab,-16'h00b8,-16'h0028,-16'h001b,-16'h0129,-16'h003a,16'h0114,-16'h0073,-16'h017b,16'h00b8,16'h005f,-16'h009b,-16'h00da,-16'h0158,16'h0171,16'h0084,16'h0047,16'h0046,16'h0026,16'h0066,-16'h01a3,-16'h00e1,-16'h0072,16'h0291,16'h0047,-16'h037d,16'h0084,-16'h0004,-16'h00ad,16'h00d4,16'h015b,16'h001e,-16'h0016,16'h003c,16'h0096,-16'h01c4,16'h019e,16'h0023,-16'h0223,-16'h008c,-16'h01c1,16'h00a6,-16'h0371,-16'h0013,-16'h013d,16'h0107,-16'h006c,16'h0140,16'h0082,-16'h006d,16'h00b0,-16'h0056,16'h0188,-16'h00c5,16'h019d,16'h0010,16'h00e2,16'h0000,-16'h017a,16'h00df,-16'h009b,-16'h00a7,16'h0286,16'h01d6,-16'h000f,-16'h0093,16'h004d,16'h00c0,-16'h00a7,-16'h008a,16'h00e1,-16'h001f,-16'h00e7,16'h0026,16'h001f,-16'h0092,-16'h00d2,-16'h00ad,16'h0147,16'h006c,-16'h006c,16'h0038,16'h0024,16'h0112,-16'h0143,-16'h0112,-16'h00c8,16'h02dc,16'h00b0,-16'h02d8,16'h00e1,16'h001b,-16'h00c4,16'h00dd,16'h0143,16'h001b,16'h0041,-16'h0072,16'h00bc,-16'h0128,16'h00f6,-16'h0053,-16'h0108,-16'h000f,-16'h00dd,16'h00ee,-16'h02ee,-16'h004d,-16'h0115,-16'h0035,-16'h008f,16'h0071,16'h00a0,-16'h00a0,16'h00e6,16'h004f,16'h0148,-16'h0108,16'h0204,-16'h008c,16'h0035,16'h0043,-16'h00d5,16'h0055,-16'h004f,-16'h004d,16'h020d,16'h015d,-16'h0025,-16'h0149,16'h0093,16'h012d,-16'h00c6,-16'h00cc,16'h00bc,-16'h0014,-16'h0083,-16'h001b,-16'h0046,16'h000e,-16'h00d3,-16'h0038,16'h0138,-16'h000c,-16'h0099,16'h0044,16'h0015,16'h0161,-16'h00ae,-16'h012e,-16'h00b2,16'h0248,16'h0157,-16'h0219,-16'h0074,16'h004b,-16'h00c6,16'h00c7,16'h01c0,16'h006a,16'h003d,-16'h000e,16'h0116,-16'h00bc,16'h0132,-16'h0094,-16'h000c,16'h0009,-16'h0052,16'h0066,-16'h015f,16'h002e,-16'h00f7,-16'h00ab,16'h0088,-16'h0055,-16'h0001,16'h005d,16'h00f6,-16'h0054,16'h0213,-16'h00f6,16'h02f9,-16'h0088,-16'h005a,-16'h0044,-16'h009d,16'h004f,-16'h0066,-16'h0069,16'h00a4,16'h0173,-16'h0093,-16'h01a6,-16'h0033,16'h00d2,-16'h0043,-16'h00a2,16'h00c1,16'h002b,-16'h000b,-16'h0094,-16'h007b,16'h00f6,16'h00eb,16'h0082,16'h0051,16'h0005,-16'h0066,16'h00f6,16'h0157,-16'h00a1,16'h00ff,16'h00ba,16'h0089,16'h00a8,-16'h005b,16'h0007,-16'h0037,-16'h009f,16'h0175,-16'h0069,16'h0027,16'h000e,-16'h0086,-16'h00e4,16'h0080,16'h0100,-16'h00eb,-16'h0070,-16'h010f,16'h00a3,-16'h005d,16'h0000,-16'h005f,16'h0144,16'h00b5,-16'h0061,-16'h0040,16'h0045,-16'h0011,16'h0127,-16'h00cb,16'h0059,16'h0198,-16'h0056,-16'h0001,-16'h0005,-16'h000a,16'h000e,16'h0061,16'h0016,16'h012c,16'h0105,-16'h0083,16'h0108,16'h000c,16'h003c,16'h0077,-16'h00c0,-16'h0085,-16'h00a3,-16'h005c,-16'h0072,16'h0016,16'h0091,-16'h0014,16'h0099,16'h00cb,16'h004f,16'h006a,-16'h0036,-16'h003e,16'h0188,16'h0092,-16'h0080,16'h00ce,16'h0083,16'h009b,16'h0159,-16'h00b7,-16'h0037,-16'h000b,16'h004e,16'h00fc,-16'h001d,-16'h0003,-16'h0075,-16'h0126,-16'h00d7,16'h0084,16'h0139,-16'h0084,-16'h0068,-16'h0131,16'h009b,-16'h0043,16'h007a,-16'h0013,16'h0206,16'h0160,16'h001e,-16'h0001,16'h0091,-16'h0073,16'h012c,-16'h0088,16'h002c,16'h0174,-16'h0025,16'h0057,-16'h0075,-16'h002c,16'h000c,16'h00b9,-16'h002d,16'h00b0,16'h00ab,-16'h0083,16'h012d,16'h0043,16'h003d,16'h0080,-16'h00a3,-16'h0081,-16'h00fc,-16'h0060,-16'h00a4,-16'h007f,16'h00a8,-16'h0051,16'h007b,16'h00b1,16'h0019,16'h00c2,-16'h002c,-16'h00b5,16'h017b,16'h003a,-16'h0126,16'h012d,16'h00c9,16'h0050,16'h0211,-16'h00ff,-16'h0022,-16'h007f,16'h006c,16'h00b1,-16'h003e,-16'h0082,-16'h0079,-16'h00f8,-16'h00f8,16'h007e,16'h00f7,-16'h009d,-16'h004a,-16'h0112,16'h0060,-16'h0014,16'h0055,16'h000e,16'h02ba,16'h0193,16'h00d3,-16'h0022,16'h006a,16'h000c,16'h011e,-16'h00ce,-16'h0004,16'h00ff,-16'h0061,16'h0088,-16'h00c3,16'h001f,16'h0024,16'h00c2,-16'h0041,16'h00c6,16'h00ad,-16'h012d,16'h013b,-16'h0022,16'h003f,16'h00e1,-16'h0082,-16'h0031,-16'h0131,-16'h0037,-16'h0105,-16'h0058,16'h00d1,-16'h002d,16'h0071,16'h010e,16'h0012,16'h00e8,-16'h0068,-16'h00a0,16'h01a6,16'h003d,-16'h0128,16'h00fa,-16'h0028,16'h0063,16'h0176,-16'h0136,-16'h00ad,16'h0067,16'h00a0,16'h004a,16'h0027,-16'h00bc,-16'h0033,-16'h013b,-16'h0057,16'h0013,16'h00a1,16'h000d,16'h0053,-16'h019d,16'h004e,16'h0000,16'h0000,-16'h0004,16'h0259,16'h0165,16'h0028,-16'h00be,16'h0103,16'h001e,16'h00f1,-16'h0095,-16'h006f,16'h013c,-16'h0027,16'h0037,-16'h0137,16'h0026,-16'h0038,16'h007e,-16'h005e,16'h004c,16'h002d,-16'h0124,16'h0135,16'h0001,-16'h0013,16'h0174,-16'h00bd,-16'h0034,-16'h00fd,-16'h008a,-16'h00eb,16'h0018,16'h0030,16'h0070,16'h003f,16'h010f,16'h0067,16'h007e,-16'h0040,-16'h0022,16'h0214,-16'h003f,-16'h007e,16'h00f9,-16'h00b9,-16'h0004,16'h0238,-16'h0132,-16'h0150,16'h0050,16'h001e,-16'h002c,-16'h002e,-16'h0119,-16'h0026,-16'h01a1,16'h0054,-16'h0065,16'h0116,16'h0027,16'h008d,-16'h0183,16'h0063,16'h0024,-16'h0009,16'h005f,16'h025e,16'h00fe,16'h006b,-16'h00ce,16'h016a,-16'h00e1,16'h0106,-16'h0001,-16'h006a,16'h00e4,-16'h0105,16'h0031,-16'h018e,16'h0092,-16'h00a7,16'h00a1,16'h0023,-16'h006b,16'h0020,-16'h0160,16'h0086,-16'h005e,-16'h0056,16'h006f,-16'h00de,-16'h0080,-16'h01ca,-16'h0141,-16'h005b,16'h003c,16'h00b4,16'h003c,16'h0070,16'h0054,16'h0071,16'h0058,-16'h0063,16'h0088,16'h0184,16'h002c,-16'h0035,16'h0062,-16'h01a7,16'h0028,16'h0125,-16'h0112,-16'h0255,16'h00b3,16'h005d,16'h0039,16'h0002,-16'h01e2,16'h0000,-16'h0124,16'h00b2,-16'h0122,16'h0046,16'h0006,16'h0136,-16'h0079,16'h00ee,-16'h002b,-16'h0064,16'h0014,16'h01ab,16'h00ad,16'h0013,-16'h00db,16'h017f,-16'h0167,-16'h0017,16'h0062,-16'h001a,16'h0177,-16'h00c6,-16'h0013,-16'h01b2,16'h00f0,-16'h0119,16'h0068,16'h0030,-16'h00ac,-16'h005b,-16'h00d8,16'h00c8,-16'h0008,-16'h00bb,16'h0025,-16'h0079,16'h004e,-16'h014e,-16'h022d,16'h005f,16'h0045,16'h010d,16'h0039,-16'h002a,16'h0036,16'h00ba,16'h00b5,-16'h014f,16'h00b6,16'h01b3,-16'h0002,-16'h0052,16'h00c3,-16'h0204,16'h00c9,16'h00ba,-16'h003a,-16'h02d2,16'h00ee,16'h00ff,16'h005a,-16'h0021,-16'h01c9,-16'h003d,-16'h003a,16'h01bf,-16'h00ac,16'h008b,16'h0067,16'h00ec,-16'h011c,16'h0069,16'h0051,-16'h01ac,16'h008c,16'h0124,16'h002f,16'h0031,-16'h00cb,16'h0118,-16'h022a,16'h0030,16'h0003,-16'h00b7,16'h0186,16'h0068,-16'h006f,-16'h012c,16'h002c,-16'h00ee,-16'h0015,-16'h0025,-16'h00f6,-16'h002a,16'h000b,16'h00db,-16'h0003,-16'h0040,-16'h0021,-16'h00fa,-16'h0024,-16'h01aa,-16'h028b,16'h0018,16'h00dd,16'h01a5,16'h00b4,-16'h00f8,16'h0014,16'h00bb,16'h013b,-16'h0204,16'h0092,16'h0189,16'h0068,16'h0013,16'h0034,-16'h0308,16'h0079,16'h0096,16'h005f,-16'h0369,16'h003e,16'h0118,16'h008c,-16'h008c,-16'h00c4,16'h0068,-16'h0003,16'h00c6,16'h0011,16'h00ae,16'h0058,16'h00c2,-16'h00a4,-16'h0048,-16'h009f,-16'h01c8,16'h006b,16'h00ef,16'h0022,16'h0015,-16'h004e,16'h00e7,-16'h01ae,-16'h001e,16'h0053,-16'h010c,16'h0190,16'h00f7,-16'h00a0,-16'h0095,-16'h008d,-16'h00a2,16'h0084,-16'h0050,-16'h00ef,-16'h003d,16'h007e,16'h00e1,16'h006d,-16'h001a,-16'h0095,-16'h0156,16'h00b1,-16'h018e,-16'h02c2,16'h0028,16'h00ab,16'h01b8,16'h000a,-16'h009f,-16'h0026,16'h005c,16'h010f,-16'h02d8,16'h0106,16'h00ec,16'h00de,16'h0031,16'h0004,-16'h02a3,16'h010e,16'h0062,16'h00e0,-16'h0477,-16'h000e,16'h00f4,16'h0048,-16'h018d,-16'h008b,16'h0034,16'h0017,16'h00f1,16'h001f,16'h00bc,16'h0086,-16'h0018,16'h0030,-16'h0022,-16'h0055,-16'h0132,-16'h0031,-16'h0009,-16'h000c,-16'h002f,-16'h0033,16'h0077,16'h0029,-16'h00d5,16'h001f,-16'h0115,16'h01ca,16'h00ad,-16'h0153,-16'h0073,-16'h00d8,-16'h005a,16'h0082,-16'h0028,-16'h00b2,16'h002c,16'h00ae,16'h0128,16'h0094,16'h0016,-16'h0131,-16'h016e,16'h00b8,-16'h01c8,-16'h0308,16'h0102,16'h011f,16'h0127,-16'h0006,-16'h004c,16'h0012,-16'h0050,16'h011e,-16'h0397,16'h0116,16'h00b1,16'h00d7,16'h0044,-16'h00a6,-16'h02f7,16'h0182,16'h00ee,16'h00d2,-16'h0596,-16'h0037,16'h0103,-16'h0012,-16'h0235,-16'h00f6,-16'h0036,-16'h000e,16'h0088,16'h00a5,16'h00dc,16'h0013,-16'h0154,16'h00e6,-16'h0056,-16'h004b,-16'h00cd,-16'h0083,-16'h00a5,-16'h0024,-16'h0090,16'h001a,-16'h0068,16'h0052,-16'h00ac,-16'h0148,-16'h0028,16'h01c6,16'h0030,-16'h0077,-16'h0090,-16'h0082,-16'h008c,16'h005a,16'h0024,16'h000d,-16'h003e,16'h010a,16'h00fe,16'h00c8,-16'h0044,-16'h00d4,-16'h0117,16'h0024,-16'h017b,-16'h0270,16'h00a2,16'h0192,16'h011e,-16'h0064,-16'h001b,-16'h0021,-16'h002e,16'h0161,-16'h0345,16'h016f,16'h00ff,16'h00a2,16'h0009,-16'h002b,-16'h02dc,16'h00f7,16'h0089,16'h0177,-16'h0615,-16'h00f5,16'h0061,16'h001d,-16'h0189,-16'h00f1,16'h008e,-16'h00eb,16'h0078,16'h0010,16'h0118,16'h006e,-16'h0148,16'h00a0,-16'h00b0,-16'h00bf,16'h0036,-16'h00aa,-16'h00e3,-16'h0120,16'h0001,16'h004f,16'h0058,16'h0008,-16'h00c5,-16'h0261,-16'h0045,16'h0136,-16'h0011,-16'h0021,-16'h0057,16'h001a,-16'h0005,16'h00ac,16'h0090,16'h003a,-16'h0017,16'h00ff,16'h00fe,16'h0060,-16'h000a,-16'h0073,-16'h003b,16'h0121,-16'h0124,-16'h02a1,16'h0100,16'h00ee,16'h00d2,16'h0008,-16'h000f,-16'h0048,-16'h00ac,16'h0127,-16'h0372,16'h011c,16'h0073,16'h00c9,-16'h0066,16'h0057,-16'h023c,16'h0125,-16'h0085,16'h0117,-16'h06b0,-16'h0047,16'h0052,16'h0040,-16'h004e,-16'h013e,16'h007c,-16'h00b4,16'h0045,16'h006e,16'h0042,16'h003e,-16'h00c5,16'h0063,-16'h0047,-16'h00b9,16'h0135,-16'h0090,-16'h00a9,-16'h01b9,16'h0094,16'h00bc,16'h0042,-16'h00c6,-16'h0078,-16'h016f,-16'h0080,16'h00d0,-16'h0008,16'h00b2,-16'h0096,16'h003d,-16'h0029,16'h0010,16'h0026,-16'h002d,-16'h00cf,16'h0082,16'h008d,-16'h0001,-16'h0079,-16'h00d5,-16'h0031,16'h00b2,-16'h00c3,-16'h02b0,16'h008f,16'h0117,16'h0025,-16'h004e,-16'h0042,16'h0009,-16'h0127,16'h00af,-16'h02f6,16'h0121,16'h00db,16'h009a,-16'h014c,16'h0132,-16'h024d,16'h010d,-16'h016d,16'h010a,-16'h06f2,-16'h004c,-16'h0002,16'h00c4,16'h00dc,-16'h0140,16'h0094,16'h0094,16'h0056,16'h0127,16'h0033,16'h0098,-16'h007c,-16'h0001,-16'h0009,-16'h0093,16'h0180,-16'h009a,-16'h00b6,-16'h0149,16'h0068,-16'h0092,-16'h0030,-16'h00c3,-16'h00ed,-16'h0175,-16'h0032,16'h01a0,16'h0007,16'h007d,-16'h0024,-16'h0051,16'h000c,-16'h005a,16'h00a9,-16'h0030,-16'h0050,-16'h003e,16'h0085,16'h0038,-16'h0027,-16'h00b8,16'h0035,16'h0037,-16'h00fb,-16'h038b,16'h0041,16'h0125,-16'h003b,-16'h0074,-16'h00f3,16'h0083,-16'h0097,16'h00f5,-16'h0225,16'h004e,16'h009f,16'h010c,-16'h014f,16'h0171,-16'h0193,16'h011b,-16'h0028,16'h008e,-16'h05fa,-16'h0025,16'h0083,16'h009b,16'h00cd,-16'h01f5,16'h001a,16'h00bc,16'h004a,16'h009c,-16'h001d,16'h0008,16'h00e6,-16'h0143,-16'h0013,-16'h0126,16'h0111,-16'h00a9,-16'h0169,-16'h00c6,16'h00db,-16'h009c,-16'h0049,-16'h0049,-16'h0104,-16'h002d,-16'h000b,16'h01ce,-16'h0058,-16'h002b,-16'h001b,-16'h001f,-16'h000e,-16'h0138,16'h004a,-16'h0044,16'h0042,-16'h0106,16'h0088,16'h008e,16'h0034,-16'h0061,16'h002a,-16'h0084,-16'h00ee,-16'h04ea,-16'h006c,16'h00e0,-16'h00ef,-16'h00ee,-16'h0087,16'h00ce,-16'h004c,16'h0108,-16'h0120,-16'h000d,16'h00c3,16'h014a,-16'h00c7,16'h0130,-16'h0208,16'h0135,16'h002f,16'h00bd,-16'h05fc,-16'h004a,-16'h000f,-16'h0014,16'h0143,-16'h01d3,-16'h002b,16'h003a,16'h0094,16'h0063,-16'h0039,16'h0086,16'h00d7,-16'h00df,16'h0089,-16'h0146,16'h00e0,-16'h0016,-16'h0168,-16'h000e,16'h00f5,-16'h00f3,-16'h0002,16'h001e,-16'h00f9,16'h0090,16'h0050,16'h0237,-16'h0020,16'h004d,16'h012a,-16'h0064,16'h0032,-16'h0190,16'h0021,-16'h007a,16'h006e,-16'h010e,16'h00af,16'h0035,-16'h0012,-16'h00cb,16'h00c3,-16'h0154,-16'h0042,-16'h0488,-16'h00a2,16'h0044,-16'h0104,-16'h0079,-16'h0087,16'h0095,16'h005f,16'h01a6,-16'h0043,16'h0085,16'h0112,16'h0108,-16'h0017,16'h00ba,-16'h0228,16'h0119,-16'h001e,16'h0053,-16'h05d6,-16'h0095,-16'h001a,16'h004a,16'h0050,-16'h0283,-16'h006c,-16'h002c,16'h001a,16'h001a,-16'h0035,16'h0091,16'h0184,-16'h005a,16'h014f,-16'h019e,-16'h0022,-16'h007f,-16'h013d,-16'h0012,16'h0084,-16'h00e1,-16'h0056,16'h0165,-16'h0114,16'h013c,16'h006a,16'h025e,16'h0025,-16'h0073,16'h01b5,-16'h0079,16'h0068,-16'h0144,-16'h003a,-16'h00b9,16'h00e2,-16'h012d,16'h0158,16'h0102,-16'h0026,-16'h0191,16'h0006,-16'h00f8,-16'h0078,-16'h042e,-16'h0041,-16'h006c,-16'h00f1,-16'h0040,-16'h0030,16'h0059,16'h003a,16'h0220,-16'h0001,16'h0000,16'h014e,16'h0189,-16'h004a,16'h004e,-16'h02f1,16'h0048,16'h0088,-16'h0057,-16'h0585,16'h003b,16'h0017,-16'h005e,-16'h0077,-16'h022f,-16'h0033,-16'h0037,16'h0037,16'h0000,-16'h0045,16'h00ae,16'h00b5,-16'h003d,16'h0137,-16'h012a,-16'h01c6,16'h0022,-16'h0133,16'h006f,16'h0154,-16'h00fb,16'h0055,16'h014c,-16'h016c,16'h0156,16'h00ff,16'h0236,16'h0077,16'h002b,16'h01d3,-16'h0078,16'h009c,-16'h0221,16'h002d,-16'h012c,16'h00c4,-16'h0129,16'h00bb,16'h00b6,-16'h0005,-16'h00ea,16'h0083,-16'h0020,-16'h0069,-16'h03d4,-16'h002f,-16'h00ca,-16'h002a,-16'h0057,16'h008a,16'h0049,16'h0033,16'h0206,-16'h00d2,16'h0010,16'h00ad,16'h0109,16'h0053,16'h0077,-16'h02ed,16'h001d,-16'h003f,16'h0030,-16'h057a,16'h00aa,16'h0021,16'h0006,16'h001f,-16'h021a,-16'h0029,-16'h004f,16'h005e,-16'h0033,-16'h00d1,16'h00e7,16'h00c5,-16'h00ec,16'h00aa,-16'h0101,-16'h0118,16'h004d,-16'h01cd,16'h0026,16'h0145,-16'h00e6,16'h00c2,16'h01ab,-16'h01a4,-16'h0064,16'h00b9,16'h01f4,-16'h001d,16'h00eb,16'h0197,-16'h004b,16'h00ac,-16'h02ba,-16'h003d,-16'h00b9,16'h0063,-16'h0169,16'h012d,16'h00c6,-16'h005c,-16'h0133,16'h008d,16'h00ac,-16'h004a,-16'h0386,-16'h001f,-16'h00fa,16'h000f,-16'h006e,16'h00e3,16'h0027,16'h00b4,16'h01e0,-16'h007f,16'h003d,16'h00f0,16'h00b5,16'h00a6,16'h006f,-16'h01f6,-16'h0068,-16'h0076,16'h0029,-16'h0583,16'h00ea,-16'h00b4,-16'h0118,16'h006e,-16'h015f,-16'h00c0,-16'h0108,16'h00a3,16'h003d,-16'h00fe,16'h0122,16'h0031,-16'h0053,16'h00cc,-16'h0171,-16'h00bd,16'h00c8,-16'h0188,16'h0011,16'h0117,16'h0023,16'h012a,16'h0007,-16'h010c,-16'h014f,16'h00b6,16'h01c9,-16'h003d,16'h014e,16'h00f5,-16'h0001,16'h007a,-16'h02e3,-16'h0030,-16'h007c,-16'h0049,-16'h0141,16'h0147,16'h0086,16'h0044,-16'h016f,16'h0007,16'h0082,16'h003d,-16'h0300,16'h005c,-16'h0126,16'h001e,-16'h001f,16'h012e,16'h0065,-16'h0077,16'h017d,-16'h000c,-16'h0016,16'h0120,16'h00a3,16'h0015,16'h00c8,-16'h0191,16'h0020,-16'h00af,16'h00e6,-16'h045d,16'h010a,16'h0000,-16'h00bd,16'h00f1,-16'h0116,-16'h00ce,-16'h0109,16'h0181,-16'h001c,-16'h0121,16'h00e9,16'h008a,16'h004b,-16'h0005,-16'h011d,-16'h0086,16'h0052,-16'h01a7,-16'h003f,16'h00c2,16'h0102,16'h0149,-16'h009d,-16'h0026,-16'h0297,16'h00ac,16'h019f,16'h0028,16'h01ba,16'h00f9,-16'h003d,16'h0035,-16'h0266,16'h0033,-16'h0100,-16'h00ea,-16'h0133,16'h0187,16'h0096,-16'h0090,-16'h014b,-16'h0082,16'h00b7,16'h00a6,-16'h029d,16'h000a,-16'h0132,-16'h006f,16'h0006,16'h016b,16'h00f6,-16'h0112,16'h0159,-16'h004c,-16'h001a,16'h0099,16'h00c0,16'h003b,16'h0045,-16'h0195,-16'h006a,16'h0001,16'h0040,-16'h041b,16'h00d6,16'h001c,-16'h0149,16'h00fc,-16'h016a,-16'h00d6,-16'h00d3,16'h0245,16'h0013,-16'h01e2,16'h01a2,-16'h003b,16'h005a,-16'h02d1,-16'h0123,-16'h0032,16'h0093,-16'h0107,-16'h00ea,16'h00cc,16'h017d,16'h01aa,-16'h0095,16'h0072,-16'h01cb,16'h00d2,16'h01f2,16'h0059,16'h0160,16'h0097,-16'h003b,16'h0063,-16'h0206,16'h005b,-16'h00bf,-16'h00be,-16'h01d6,16'h01ae,16'h00c0,-16'h00cd,-16'h00f8,-16'h0004,16'h009b,16'h0125,-16'h0252,16'h000b,-16'h0267,16'h005e,16'h0072,16'h00cd,16'h00d7,-16'h0116,16'h021b,16'h0098,-16'h0007,16'h00b5,16'h00cf,16'h0049,16'h0055,-16'h012c,-16'h003f,16'h008c,16'h00d6,-16'h03ef,16'h00cc,16'h0005,-16'h00b3,16'h003e,-16'h00ed,-16'h0189,-16'h00a0,16'h021c,16'h0017,-16'h025d,16'h01ea,-16'h00b0,-16'h001c,-16'h062e,-16'h00fa,16'h000f,16'h0074,-16'h00d4,-16'h0198,16'h0087,16'h01c8,16'h019a,16'h0014,16'h002b,16'h000f,16'h00a6,16'h01cf,16'h0066,16'h01a9,-16'h0018,-16'h007e,-16'h0008,-16'h0160,16'h0025,-16'h0113,-16'h010a,-16'h0121,16'h0177,16'h00d3,-16'h012e,-16'h011e,16'h0044,16'h006a,16'h0145,-16'h0193,-16'h0034,-16'h0365,16'h0078,16'h00de,16'h0098,16'h0053,-16'h01f6,16'h01f2,16'h015f,-16'h000c,16'h00a9,16'h00dc,-16'h003a,-16'h0043,-16'h01a7,16'h008a,16'h013a,16'h00af,-16'h0338,16'h0065,16'h00e3,-16'h00a8,-16'h00b1,-16'h00c1,-16'h0101,-16'h0095,16'h01cb,16'h0011,-16'h0224,16'h01d8,-16'h004d,-16'h011b,-16'h0599,-16'h0172,-16'h000b,16'h002e,-16'h00a1,-16'h00b9,16'h00ca,16'h0231,16'h0147,-16'h0020,16'h004a,16'h00bb,16'h0089,16'h01ba,16'h0078,16'h0131,-16'h003e,-16'h003c,16'h0020,-16'h0140,16'h0001,-16'h00f4,-16'h0111,-16'h000b,16'h01de,16'h0041,-16'h0190,-16'h00cc,16'h003c,-16'h00db,16'h0165,-16'h00d4,16'h0017,-16'h0411,16'h0028,16'h00b3,16'h0039,-16'h0049,-16'h0187,16'h010d,16'h0139,16'h0023,16'h0057,-16'h0001,16'h0037,-16'h00e1,-16'h0107,16'h00b7,16'h0166,16'h0128,-16'h0372,16'h0087,16'h0152,-16'h014c,-16'h0117,-16'h0098,16'h0027,-16'h00d7,16'h00d3,16'h0079,-16'h0285,16'h01ed,16'h0058,-16'h020d,-16'h0348,-16'h0196,16'h005d,-16'h0070,-16'h00bd,-16'h00e3,16'h010e,16'h01d2,16'h0193,16'h007d,-16'h000b,16'h0089,16'h0090,16'h0228,-16'h00b7,16'h01ad,-16'h005d,16'h0028,16'h00b7,-16'h016e,16'h0080,-16'h013c,-16'h00ea,16'h0139,16'h0283,-16'h0084,-16'h01d3,-16'h00f9,16'h006d,-16'h018c,16'h0076,-16'h0089,-16'h0004,-16'h0273,16'h00a0,16'h00ec,16'h004b,-16'h015f,-16'h012c,16'h009f,16'h0198,16'h0067,16'h0082,-16'h0034,16'h008c,-16'h0170,-16'h00b2,16'h001a,16'h02af,16'h011b,-16'h0344,16'h000c,16'h0083,-16'h00e2,16'h0024,-16'h0049,-16'h002b,-16'h0097,16'h00cb,16'h00ad,-16'h022b,16'h021e,16'h004f,-16'h0204,-16'h0171,-16'h01b9,16'h00b7,-16'h0291,-16'h0053,-16'h0136,16'h0058,16'h00e6,16'h019f,16'h003f,-16'h005d,16'h0115,16'h00a4,16'h0270,-16'h01c9,16'h013b,-16'h0080,-16'h0019,16'h002f,-16'h014c,16'h0061,-16'h00a2,-16'h00ff,16'h0203,16'h0191,-16'h00b1,-16'h022f,-16'h00a7,16'h00ad,-16'h015a,-16'h0122,-16'h00be,16'h0005,-16'h0139,16'h0105,16'h0084,16'h0060,-16'h0159,-16'h0087,16'h01ad,16'h005f,16'h0057,16'h00b7,-16'h0016,16'h012f,-16'h0121,-16'h00cf,-16'h0048,16'h03ba,16'h0127,-16'h02bb,16'h007a,-16'h0031,-16'h005a,16'h0017,16'h0014,16'h0043,-16'h001a,16'h00b2,16'h00c6,-16'h01d6,16'h0175,16'h0014,-16'h01d7,-16'h0081,-16'h0138,16'h00a7,-16'h038a,16'h0018,-16'h00b3,16'h0039,16'h00da,16'h00b5,16'h00b1,-16'h006c,16'h00dc,16'h0072,16'h02b5,-16'h01ec,16'h0212,-16'h0048,-16'h0060,16'h0058,-16'h010f,16'h00e0,-16'h004e,-16'h00c3,16'h018e,16'h019e,-16'h0096,-16'h0143,-16'h0017,16'h01a4,-16'h0108,-16'h0152,-16'h0039,-16'h00fd,-16'h001e,-16'h0008,16'h000b,16'h0035,-16'h0112,-16'h002f,16'h0175,-16'h002a,-16'h0021,16'h009a,16'h0022,16'h01b1,-16'h0111,-16'h0062,-16'h008b,16'h033e,16'h0095,-16'h0247,16'h0060,-16'h0015,-16'h008f,-16'h0013,16'h002b,16'h0001,16'h0051,16'h0083,16'h0183,-16'h0185,16'h0145,-16'h008b,-16'h00f7,-16'h000c,-16'h0086,16'h0046,-16'h0275,-16'h0014,-16'h00ff,-16'h0092,16'h00b0,16'h00a5,16'h00b2,-16'h0074,16'h0049,16'h001a,16'h02f7,-16'h018c,16'h0281,-16'h0074,-16'h00ec,16'h000e,-16'h00f0,16'h0083,16'h0021,-16'h002c,16'h019d,16'h0146,-16'h0083,-16'h0119,16'h000a,16'h017f,-16'h0058,-16'h0149,-16'h00a6,-16'h0043,16'h002c,-16'h003c,16'h0025,16'h005e,-16'h00e1,-16'h0018,16'h0139,-16'h003f,-16'h0120,16'h0048,-16'h0031,16'h01bf,-16'h00cd,-16'h007e,16'h0012,16'h029a,16'h00c1,-16'h01bb,-16'h001d,16'h0052,-16'h004e,16'h0036,16'h01a1,16'h0085,-16'h0017,16'h001f,16'h014c,-16'h00d2,16'h0172,-16'h0054,-16'h0035,16'h0002,-16'h0039,16'h0070,-16'h017f,16'h0001,-16'h004e,-16'h0120,16'h00ac,-16'h0065,16'h0005,16'h0046,16'h0066,-16'h0035,16'h0279,-16'h015b,16'h027d,-16'h0074,-16'h00e8,-16'h0011,-16'h0065,16'h0034,16'h0028,-16'h008e,16'h00e7,16'h00bb,-16'h00dd,-16'h01ba,16'h0037,16'h0171,-16'h009f,-16'h0124,-16'h0047,-16'h000f,-16'h0015,-16'h00b4,-16'h0065,16'h006c,16'h0054,16'h0030,16'h0000,-16'h003c,16'h0002,16'h003a,16'h00a0,-16'h000d,16'h0060,16'h0051,-16'h0010,16'h0068,16'h0047,-16'h0050,-16'h0023,-16'h003f,16'h00a0,-16'h002d,-16'h0043,-16'h004b,-16'h004b,-16'h0092,-16'h0029,16'h0031,-16'h0055,-16'h0018,-16'h005c,16'h0009,16'h0000,-16'h0021,-16'h0004,16'h0076,16'h0095,-16'h0012,-16'h0015,16'h0097,-16'h0076,16'h00b9,-16'h0050,-16'h0005,16'h00c8,16'h0048,16'h0000,-16'h0005,-16'h0032,16'h000e,16'h0031,-16'h0034,16'h0060,16'h009d,-16'h00b4,16'h009f,16'h0010,16'h0093,16'h0089,-16'h0003,-16'h004f,-16'h0060,-16'h005d,-16'h0033,-16'h0045,16'h004b,-16'h0027,16'h0046,16'h007f,16'h002c,16'h0022,-16'h0024,16'h0000,16'h0083,16'h0051,-16'h0048,16'h010e,16'h0039,-16'h0012,16'h0102,-16'h001a,-16'h0052,-16'h0018,-16'h0044,16'h0062,-16'h0014,16'h000a,-16'h003a,-16'h0094,-16'h00a2,16'h0026,16'h00eb,-16'h0038,-16'h0012,-16'h00b6,16'h0008,-16'h000e,-16'h0079,-16'h009e,16'h0193,16'h00d3,-16'h001f,-16'h006f,16'h0009,-16'h0006,16'h00d8,-16'h0099,16'h0053,16'h0064,-16'h002e,16'h0022,-16'h006b,16'h0018,16'h0016,16'h002e,16'h003f,16'h00d8,16'h0022,-16'h00cf,16'h00ce,-16'h0091,16'h001f,16'h008b,-16'h0034,-16'h00a9,-16'h0056,-16'h0049,-16'h0065,-16'h0065,16'h0046,16'h0024,16'h0076,16'h0196,16'h001a,16'h0077,-16'h0017,-16'h0007,16'h00f3,16'h009a,-16'h00a3,16'h0163,-16'h0009,16'h002a,16'h014a,-16'h0002,-16'h0066,-16'h0026,16'h002b,16'h00a7,-16'h0099,-16'h0049,-16'h000a,-16'h0061,-16'h001c,16'h0052,16'h00bd,-16'h0020,16'h0053,-16'h00b4,16'h0034,16'h0006,-16'h006f,-16'h0040,16'h021b,16'h00cb,16'h0030,16'h000f,16'h00cc,-16'h0017,16'h0094,-16'h0005,16'h001a,16'h0105,-16'h0071,16'h000d,-16'h0033,-16'h0027,16'h0059,16'h0047,-16'h004b,16'h0054,16'h002a,-16'h0065,16'h0068,-16'h0064,-16'h0044,16'h0085,-16'h002a,-16'h0086,-16'h00d3,-16'h0032,-16'h0119,-16'h000f,-16'h002d,-16'h001e,16'h0013,16'h01b3,-16'h006d,16'h0095,-16'h0038,-16'h0070,16'h0163,16'h0006,-16'h0043,16'h01a5,-16'h0090,16'h003b,16'h011d,-16'h0094,-16'h00c1,16'h002b,16'h0041,16'h0039,-16'h004d,-16'h0065,-16'h0085,-16'h0135,-16'h0009,-16'h0026,16'h0160,-16'h004b,16'h001a,-16'h00b5,-16'h0060,-16'h0011,-16'h0068,16'h0015,16'h021f,16'h00fe,-16'h0018,-16'h006f,16'h00fe,-16'h0057,16'h013f,16'h001f,-16'h0027,16'h00af,-16'h002b,16'h0031,-16'h0063,16'h0026,16'h0003,16'h0046,-16'h007c,16'h003e,16'h004e,-16'h0082,16'h00d5,-16'h0011,-16'h00ab,16'h0053,-16'h00b7,-16'h0042,-16'h00cb,-16'h0026,-16'h00ff,-16'h0043,16'h0038,16'h0048,-16'h0010,16'h011b,16'h0037,16'h006e,-16'h0053,16'h0082,16'h0165,16'h000b,-16'h00e7,16'h015d,-16'h0130,16'h000d,16'h0167,-16'h0083,-16'h00b3,16'h0052,-16'h001a,16'h0045,-16'h00db,-16'h005f,-16'h004f,-16'h00e1,16'h002e,-16'h0057,16'h0123,-16'h005b,16'h00a7,-16'h007e,-16'h0009,16'h003e,-16'h00a1,16'h0074,16'h024f,16'h007e,16'h005b,-16'h00e0,16'h0173,-16'h000b,16'h0129,-16'h000c,16'h0014,16'h0049,-16'h0070,16'h0099,-16'h0134,16'h0065,-16'h0072,16'h0077,16'h000f,-16'h0064,-16'h0015,-16'h00d6,16'h008b,-16'h0054,-16'h0082,16'h000a,-16'h00cc,-16'h0097,-16'h016c,-16'h00de,-16'h00b8,16'h0047,16'h0083,16'h0067,-16'h0017,16'h019b,16'h0007,16'h0089,-16'h00ab,16'h00b5,16'h013a,-16'h002c,-16'h0038,16'h0115,-16'h0139,-16'h000e,16'h0142,-16'h0055,-16'h0174,16'h0120,16'h005b,16'h009d,-16'h00fe,-16'h0127,-16'h0042,-16'h005d,16'h005b,-16'h00d3,16'h00ef,-16'h002d,16'h00c3,-16'h00e8,16'h0092,16'h000b,-16'h016d,16'h005c,16'h0266,16'h0067,-16'h001f,-16'h00b1,16'h00c5,-16'h006d,16'h00b3,-16'h000e,-16'h0050,16'h006e,-16'h0069,16'h0051,-16'h011d,16'h005b,-16'h00b1,16'h00aa,-16'h0003,-16'h0091,-16'h0009,-16'h0083,16'h005e,-16'h0008,-16'h003d,-16'h0027,-16'h0175,-16'h0024,-16'h0137,-16'h0122,-16'h0019,16'h006a,16'h00de,16'h0035,-16'h0056,16'h00c5,16'h00d3,16'h0055,-16'h00af,16'h0111,16'h00f2,-16'h008a,16'h0004,16'h0131,-16'h01db,16'h0041,16'h0165,-16'h0089,-16'h0222,16'h00e9,16'h009b,16'h0084,-16'h0124,-16'h00e1,16'h0034,16'h0019,16'h00a8,-16'h0096,16'h012f,-16'h0006,16'h014b,-16'h009b,-16'h0019,16'h0077,-16'h021e,-16'h0013,16'h0165,16'h0029,16'h0010,-16'h0031,16'h0070,-16'h0085,16'h00c2,16'h002e,-16'h0049,16'h0110,16'h0083,16'h0027,-16'h0152,16'h004d,-16'h00ba,16'h008c,-16'h0088,-16'h0125,16'h0050,-16'h004a,16'h002f,16'h0040,-16'h00b1,-16'h002e,-16'h019b,16'h0087,-16'h01be,-16'h01da,16'h0025,16'h00e5,16'h01b2,16'h0040,-16'h004e,16'h0057,16'h00e7,16'h0038,-16'h0144,16'h00c8,16'h00fc,-16'h0049,16'h0029,16'h004d,-16'h0218,16'h0033,16'h0119,16'h005d,-16'h0299,16'h007b,16'h00b6,16'h00f7,-16'h0101,-16'h00b2,16'h002d,16'h002a,16'h00a8,-16'h003f,16'h0124,-16'h0013,16'h00d7,-16'h00be,16'h0026,-16'h0007,-16'h016b,-16'h0021,-16'h0027,16'h0014,16'h000d,-16'h0068,16'h0056,-16'h0044,16'h0019,-16'h0027,-16'h00bb,16'h00b8,16'h010c,-16'h00c3,-16'h0059,16'h0018,-16'h0083,16'h00bc,-16'h007e,-16'h0135,-16'h0021,-16'h0033,16'h008c,16'h0064,-16'h0001,-16'h0083,-16'h01c1,16'h009d,-16'h01d5,-16'h01b4,-16'h0026,16'h00aa,16'h0173,16'h0067,-16'h0054,16'h009a,16'h0074,16'h0038,-16'h01c7,16'h00f7,16'h00c5,-16'h002c,16'h0058,16'h0015,-16'h01da,16'h0114,16'h012a,16'h00d4,-16'h0262,-16'h0047,16'h00c1,16'h00d3,-16'h0258,16'h001f,16'h0072,16'h0091,16'h00ad,16'h0025,16'h010d,-16'h0032,-16'h00ac,-16'h0001,-16'h00a5,-16'h001c,-16'h014e,-16'h00b1,-16'h008e,16'h0031,-16'h0022,-16'h0049,-16'h003a,16'h0073,-16'h00bc,-16'h008e,-16'h00bd,16'h00b8,16'h0085,-16'h00cc,16'h0000,-16'h001c,-16'h00c7,16'h00e3,16'h0061,-16'h008d,-16'h0081,16'h0022,16'h009c,16'h006e,16'h0017,-16'h009e,-16'h017b,16'h0064,-16'h018c,-16'h01a7,16'h00b1,16'h00d2,16'h00f4,16'h005b,-16'h0011,16'h00b6,-16'h0047,16'h0079,-16'h015f,16'h014d,16'h00da,-16'h000a,16'h0074,-16'h0028,-16'h023c,16'h0148,16'h00b7,16'h00fe,-16'h0303,-16'h00c4,16'h004f,16'h004f,-16'h0286,-16'h0024,16'h00e0,-16'h000c,16'h0086,16'h00c6,16'h0119,16'h0002,-16'h018f,16'h00b1,-16'h0050,-16'h00ca,-16'h0043,-16'h009c,-16'h0082,-16'h005f,-16'h0084,-16'h0096,16'h0022,16'h0035,-16'h0086,-16'h01f9,-16'h00c6,16'h0145,-16'h0015,-16'h00bb,16'h0093,-16'h00f9,-16'h0072,16'h005d,16'h0050,-16'h0082,-16'h0080,16'h0053,16'h00c4,16'h0050,-16'h0056,-16'h012f,-16'h0166,16'h00aa,-16'h0142,-16'h018e,16'h00dd,16'h013f,16'h00a3,16'h0033,-16'h00c1,-16'h0052,-16'h00b6,16'h0065,-16'h01d3,16'h015c,16'h00d4,16'h002b,16'h0085,16'h000e,-16'h01e2,16'h0167,16'h00ac,16'h017f,-16'h0323,-16'h00da,16'h0011,16'h0091,-16'h0111,-16'h0038,16'h00d1,-16'h0085,16'h006e,16'h0083,16'h00cf,16'h000e,-16'h01a9,16'h0054,-16'h0022,-16'h007c,16'h0141,-16'h00b2,-16'h0145,-16'h0167,16'h0062,16'h000e,16'h0023,-16'h005a,-16'h0081,-16'h017b,-16'h0068,16'h00fe,-16'h00ac,-16'h0012,16'h0058,-16'h0028,-16'h0047,16'h0025,16'h0049,-16'h0095,-16'h0021,16'h008e,16'h0097,16'h00ce,-16'h0064,-16'h00f9,-16'h00eb,16'h0093,-16'h0182,-16'h0187,16'h0101,16'h007e,16'h0033,16'h00cb,-16'h00ca,-16'h0035,-16'h0162,16'h007a,-16'h017a,16'h00d1,16'h003d,-16'h0003,-16'h0088,16'h006c,-16'h020a,16'h00e4,-16'h00ad,16'h0175,-16'h0334,-16'h009d,-16'h0059,16'h0049,16'h0069,-16'h005b,16'h00af,-16'h00c3,16'h00b9,16'h0093,16'h007d,16'h002e,-16'h0173,-16'h0030,-16'h0072,-16'h009a,16'h01af,-16'h0041,-16'h00fc,-16'h01a7,16'h0083,16'h0039,16'h0052,-16'h0108,-16'h00ae,-16'h0116,-16'h00ba,16'h011c,-16'h0052,-16'h005f,16'h0127,-16'h003b,-16'h004b,-16'h0075,16'h0033,-16'h0070,-16'h00cf,16'h00cb,16'h0114,16'h001c,-16'h00ae,-16'h00d1,-16'h007f,-16'h003b,-16'h0129,-16'h019e,16'h0002,16'h003f,-16'h009d,-16'h000b,-16'h008a,16'h002e,-16'h015c,16'h0085,-16'h0126,16'h00ad,16'h001f,16'h0013,-16'h00ec,16'h00fe,-16'h01f0,16'h0083,-16'h00a3,16'h00e5,-16'h0320,16'h001f,16'h0052,16'h0085,16'h00fd,-16'h0022,16'h00b5,16'h000e,16'h00ba,16'h012c,-16'h0020,16'h001d,-16'h0043,16'h0000,-16'h003a,-16'h0090,16'h01d0,-16'h0074,-16'h0181,-16'h012f,16'h00bb,-16'h00d6,-16'h001c,-16'h0065,-16'h0117,16'h001f,-16'h0058,16'h00db,-16'h002f,16'h0096,16'h0110,-16'h005e,16'h0009,-16'h011e,16'h0026,16'h0040,-16'h00e5,-16'h004a,16'h007c,16'h004c,-16'h0044,-16'h00a7,16'h0044,-16'h0056,-16'h0075,-16'h024a,-16'h0044,16'h008e,-16'h00d5,-16'h0077,-16'h0074,16'h00e2,-16'h00e0,16'h00ba,-16'h0118,16'h0007,16'h008c,16'h0088,-16'h0100,16'h0132,-16'h0163,16'h00c9,-16'h00e9,16'h003f,-16'h0392,16'h0050,16'h0062,16'h007e,16'h0136,-16'h0080,16'h0014,16'h002e,16'h00a8,16'h0141,-16'h00e4,16'h0080,16'h00ad,-16'h00a6,-16'h0008,-16'h009f,16'h016e,-16'h0023,-16'h0256,-16'h0108,16'h00cc,-16'h014c,16'h0065,-16'h001c,-16'h014a,16'h005f,-16'h007b,16'h01c5,-16'h0027,16'h0082,16'h014f,-16'h009f,-16'h0061,-16'h01c6,16'h0079,16'h0007,-16'h0033,-16'h0094,16'h00df,16'h004f,-16'h006d,-16'h0065,16'h00f5,-16'h00de,-16'h0085,-16'h02f4,-16'h0011,16'h0079,-16'h00c3,-16'h005a,-16'h0043,16'h00e6,-16'h002e,16'h00b1,-16'h0044,16'h0063,16'h007b,16'h010b,-16'h0109,16'h00ea,-16'h01bc,16'h0088,-16'h0014,16'h0055,-16'h0337,-16'h0025,-16'h002e,16'h0063,16'h0113,-16'h0119,16'h0043,16'h0050,16'h013c,16'h00b0,-16'h010d,16'h0055,16'h011d,-16'h00d2,16'h008d,-16'h0086,16'h00fb,16'h0079,-16'h01f3,-16'h0065,16'h00f1,-16'h0154,-16'h001a,16'h000b,-16'h0165,16'h018d,-16'h000e,16'h01b9,-16'h0026,-16'h001e,16'h019d,-16'h0034,-16'h000d,-16'h01ca,16'h0027,16'h0002,-16'h0003,-16'h01db,16'h0128,16'h007b,-16'h0049,-16'h0137,16'h00d8,-16'h015c,-16'h0023,-16'h03c2,-16'h002d,-16'h003a,-16'h0120,-16'h00aa,-16'h005c,16'h010d,-16'h007a,16'h0141,-16'h0004,16'h00f1,-16'h0054,16'h014d,-16'h0015,16'h005a,-16'h0183,16'h0073,16'h0021,-16'h0029,-16'h02f0,16'h0059,16'h0024,-16'h00b2,16'h0097,-16'h0141,-16'h0095,-16'h0038,16'h00df,16'h0025,-16'h0150,16'h005f,16'h00f9,-16'h00c5,16'h0047,-16'h00f5,16'h0045,16'h0052,-16'h0217,16'h0058,16'h013e,-16'h014a,16'h002c,16'h0119,-16'h014f,16'h0140,16'h002a,16'h01ee,16'h0013,-16'h004a,16'h0177,-16'h0024,16'h00e2,-16'h01f1,16'h0030,-16'h0058,16'h002a,-16'h0204,16'h017d,16'h008f,-16'h0080,-16'h0183,16'h00c8,-16'h0097,-16'h001d,-16'h0490,16'h0023,-16'h014e,-16'h012e,-16'h00af,-16'h0020,16'h00b1,16'h0054,16'h01c8,16'h0057,16'h00b3,16'h003c,16'h0118,-16'h0069,16'h007e,-16'h0145,16'h007b,16'h0042,-16'h00bf,-16'h02c3,16'h007d,16'h0014,-16'h0082,16'h002c,-16'h01d4,-16'h0055,-16'h0058,16'h0039,16'h0018,-16'h00c7,-16'h0003,16'h0069,-16'h00db,16'h00c9,-16'h009b,-16'h01d3,16'h001c,-16'h010a,16'h00c4,16'h011a,-16'h0153,16'h00a7,16'h01d3,-16'h00ec,16'h0055,16'h009e,16'h0256,16'h004d,-16'h0014,16'h0252,-16'h00b2,16'h00e8,-16'h01fb,16'h0014,16'h0022,16'h0074,-16'h01f7,16'h0165,16'h00e3,-16'h0054,-16'h0166,16'h00c8,-16'h001f,-16'h0003,-16'h052d,16'h0032,-16'h0154,-16'h007a,-16'h00c8,-16'h0023,16'h0053,-16'h000e,16'h01de,16'h003f,16'h00a7,16'h006c,16'h00e5,-16'h0041,16'h0067,-16'h0103,16'h0034,16'h0078,-16'h0072,-16'h0317,16'h0084,-16'h0007,-16'h00a4,16'h0047,-16'h0224,-16'h00e8,-16'h0087,16'h0037,16'h0014,-16'h0182,16'h0061,-16'h0007,-16'h016c,16'h0017,-16'h009f,-16'h00e2,16'h00c0,-16'h008d,16'h00d1,16'h0192,-16'h0094,16'h013c,16'h0116,-16'h01b4,-16'h0044,16'h00cc,16'h019e,16'h007b,16'h0070,16'h00de,16'h001a,16'h006e,-16'h01d4,16'h000f,-16'h005a,-16'h0084,-16'h0183,16'h0192,16'h00cc,-16'h0038,-16'h0208,16'h0093,16'h0070,16'h0073,-16'h0551,-16'h005d,-16'h00ae,16'h0073,-16'h003b,16'h0019,16'h00b2,-16'h008b,16'h01ed,16'h0066,16'h00c3,16'h012d,16'h0167,-16'h0057,16'h0056,-16'h00c9,16'h002c,-16'h0029,-16'h0052,-16'h0290,16'h0122,-16'h002e,-16'h01c4,16'h012e,-16'h024e,-16'h0141,-16'h004b,16'h0043,-16'h009a,-16'h014b,16'h00c9,16'h0045,-16'h00a2,16'h0084,-16'h00b3,-16'h0077,16'h004e,-16'h00bf,-16'h0005,16'h00e8,16'h0028,16'h0112,-16'h0003,-16'h011d,-16'h01af,16'h006d,16'h01b9,16'h002e,16'h00d8,16'h0138,16'h0020,16'h0070,-16'h01f7,16'h003f,-16'h0016,-16'h00bf,-16'h0175,16'h0172,16'h00d6,-16'h004e,-16'h017e,16'h0081,16'h0141,16'h0076,-16'h0599,-16'h0007,-16'h013b,16'h006e,-16'h0047,-16'h0018,16'h00ca,-16'h014d,16'h0263,16'h004d,16'h0077,16'h0098,16'h00f5,-16'h00e4,16'h005b,-16'h009d,-16'h006f,16'h0017,16'h002c,-16'h02fa,16'h0198,-16'h0060,-16'h0238,16'h0137,-16'h025b,-16'h0158,-16'h00f8,16'h012a,-16'h004b,-16'h00d2,16'h00d7,-16'h006f,-16'h0073,-16'h0094,-16'h006b,-16'h00b8,16'h007e,-16'h002d,-16'h002f,16'h00be,16'h00e7,16'h0187,-16'h00ec,-16'h0038,-16'h0245,16'h00be,16'h01b0,16'h0080,16'h0167,16'h00f2,16'h0014,16'h006d,-16'h01c7,16'h003d,-16'h00c9,-16'h0048,-16'h012b,16'h01ff,16'h0094,-16'h0110,-16'h0160,-16'h007c,16'h0130,16'h0109,-16'h04b7,-16'h008e,-16'h0166,16'h0016,-16'h0011,16'h0040,16'h009a,-16'h01db,16'h01c7,16'h0057,-16'h0055,16'h00e5,16'h0023,-16'h008b,16'h0060,-16'h00cc,-16'h0081,16'h0027,16'h009e,-16'h0366,16'h0123,-16'h0007,-16'h0113,16'h0150,-16'h0283,-16'h0142,-16'h0195,16'h028a,-16'h004a,-16'h0191,16'h010b,-16'h0090,-16'h0002,-16'h02db,-16'h0089,-16'h0043,16'h009a,-16'h006b,-16'h0099,16'h00d9,16'h01d0,16'h017e,-16'h006e,-16'h000e,-16'h016f,16'h0121,16'h0224,16'h0047,16'h0198,16'h002f,16'h0000,16'h0068,-16'h01cb,16'h00d2,-16'h00ab,-16'h013a,-16'h01d1,16'h0160,16'h0081,-16'h0224,-16'h018e,16'h0050,16'h00bd,16'h011d,-16'h03ee,-16'h0086,-16'h0285,-16'h002b,16'h003d,16'h00e5,16'h0015,-16'h019c,16'h0233,16'h00bb,16'h000e,16'h011d,16'h0078,-16'h0082,-16'h0031,-16'h00e3,-16'h0084,16'h015a,16'h010c,-16'h0324,16'h0034,-16'h0003,-16'h0152,16'h0000,-16'h0297,-16'h00b5,-16'h0107,16'h0239,16'h0033,-16'h01e5,16'h00f7,-16'h003a,-16'h0022,-16'h0551,-16'h005c,16'h001a,-16'h0003,-16'h007f,-16'h00b0,16'h00f9,16'h01e8,16'h0187,-16'h003a,-16'h0043,-16'h0037,16'h0101,16'h0240,-16'h0080,16'h018d,16'h008d,-16'h0095,16'h0025,-16'h017c,16'h005c,-16'h0114,-16'h00d7,-16'h0134,16'h01b3,16'h003d,-16'h01b6,-16'h0167,16'h00b5,16'h0016,16'h00ef,-16'h0384,-16'h0080,-16'h0316,16'h0087,16'h00cf,16'h011b,-16'h0039,-16'h012c,16'h0181,16'h00dd,-16'h0016,16'h010e,16'h0043,-16'h0023,-16'h00a6,-16'h00ec,16'h0028,16'h0186,16'h0167,-16'h02a9,16'h0060,16'h0066,-16'h0156,-16'h009d,-16'h0279,-16'h0050,-16'h00fa,16'h01c0,16'h0098,-16'h0240,16'h0173,-16'h006f,-16'h0100,-16'h042d,-16'h001f,-16'h0007,16'h005a,-16'h0074,-16'h0110,16'h010e,16'h01e5,16'h01e6,16'h0038,16'h0061,16'h0086,16'h0115,16'h02e9,-16'h005b,16'h01aa,16'h004c,-16'h0123,16'h0064,-16'h014d,16'h008f,-16'h00b2,-16'h00ae,16'h003a,16'h01b5,-16'h0043,-16'h0221,-16'h0134,16'h00ef,-16'h0077,16'h00d4,-16'h02ae,-16'h007e,-16'h0324,16'h00d1,16'h00a5,16'h00f9,-16'h00c3,-16'h00b0,16'h0031,16'h0131,16'h0043,16'h0034,-16'h008d,16'h00c1,-16'h0151,-16'h005d,16'h0084,16'h01f3,16'h00d5,-16'h02f8,-16'h0005,16'h005c,-16'h01ac,-16'h00eb,-16'h016e,16'h002a,-16'h0134,16'h0134,16'h00f9,-16'h021a,16'h018a,-16'h008c,-16'h01cd,-16'h023e,-16'h00b5,16'h0072,-16'h009d,-16'h0031,-16'h00e7,16'h014f,16'h0197,16'h01d1,16'h000e,16'h00a7,16'h006a,16'h016c,16'h02a2,-16'h013a,16'h014d,-16'h005d,-16'h0099,16'h0072,-16'h00ef,16'h00a0,-16'h003e,-16'h00c6,16'h0140,16'h015b,-16'h0075,-16'h024c,-16'h0109,16'h00c6,-16'h00f5,-16'h0094,-16'h0272,16'h0014,-16'h0209,16'h0100,16'h00b6,16'h0089,-16'h0182,-16'h000f,16'h00c4,16'h00aa,16'h0093,16'h0094,-16'h0035,16'h00c2,-16'h0125,-16'h0014,16'h0069,16'h031b,16'h015e,-16'h02a4,16'h003a,16'h007d,-16'h00ce,-16'h0028,-16'h0142,16'h000d,-16'h009b,16'h0130,16'h00b0,-16'h01e5,16'h0140,-16'h003a,-16'h01c0,-16'h0112,-16'h0087,16'h0083,-16'h01e7,16'h0024,-16'h017f,16'h0120,16'h01b3,16'h021f,16'h000b,16'h0080,16'h0149,16'h0109,16'h0340,-16'h0213,16'h012c,16'h0003,-16'h003d,16'h006e,-16'h00d4,16'h0041,-16'h001a,-16'h00dc,16'h0148,16'h014f,-16'h0077,-16'h01b3,-16'h000c,16'h0149,-16'h011e,-16'h0129,-16'h023f,16'h0018,-16'h010a,16'h00f5,16'h0107,16'h00cd,-16'h01ae,-16'h0019,16'h00e2,16'h001f,16'h000e,16'h00e8,-16'h00b4,16'h017a,-16'h00d7,-16'h005b,-16'h007e,16'h0306,16'h0098,-16'h022f,16'h0134,-16'h003b,-16'h009e,16'h0032,-16'h00f2,16'h0057,-16'h0026,16'h00fa,16'h015e,-16'h015f,16'h0100,-16'h0063,-16'h012f,-16'h0035,-16'h0030,16'h003d,-16'h0270,-16'h0047,-16'h00c6,-16'h001e,16'h0078,16'h019d,16'h00d1,-16'h0050,16'h00e1,16'h00a7,16'h0314,-16'h01d5,16'h01b4,-16'h0065,-16'h0100,16'h005d,-16'h0087,16'h0037,16'h0086,-16'h00b2,16'h0231,16'h00d5,-16'h00c1,-16'h0145,-16'h0012,16'h0177,-16'h00ea,-16'h00ff,-16'h0230,-16'h0067,-16'h0050,16'h0085,16'h011a,16'h00e2,-16'h0179,16'h002a,16'h0089,16'h0009,-16'h002e,16'h004b,16'h0021,16'h01e9,-16'h0086,-16'h003e,-16'h007e,16'h02fe,16'h0105,-16'h023b,16'h0031,16'h0054,-16'h0076,-16'h0037,-16'h0028,16'h00b5,16'h0035,16'h00c9,16'h0112,-16'h00c4,16'h00fa,-16'h0081,-16'h0075,-16'h0001,-16'h0029,16'h0049,-16'h01cc,-16'h000a,-16'h0072,-16'h007c,16'h00f0,16'h0001,16'h0065,16'h0013,16'h0024,-16'h0037,16'h02c6,-16'h01ce,16'h01bd,-16'h0084,-16'h0104,-16'h0070,-16'h00a5,16'h0050,-16'h0023,-16'h0028,16'h0174,16'h007c,-16'h00e4,-16'h00c9,16'h006b,16'h01e8,-16'h007f,-16'h0126,-16'h0143,-16'h004d,16'h002e,-16'h0076,16'h0017,16'h0051,-16'h008e,16'h0060,16'h009b,16'h0056,-16'h0070,16'h0039,16'h0022,16'h01d5,-16'h0009,16'h0029,16'h001c,16'h0209,16'h00dd,-16'h01bc,-16'h00c0,-16'h000f,-16'h0011,-16'h0023,16'h0078,16'h007e,16'h0047,16'h003a,16'h00a9,-16'h0080,16'h00a0,-16'h00ee,16'h0007,-16'h0017,16'h0038,-16'h005f,-16'h00d6,-16'h0019,-16'h003d,-16'h0132,16'h0057,-16'h002f,-16'h0004,16'h004f,16'h0004,-16'h0084,16'h0248,-16'h0113,16'h024d,-16'h004b,-16'h00e4,-16'h00e5,-16'h0044,16'h0074,-16'h007d,-16'h005d,16'h00e5,16'h00bf,-16'h007d,-16'h0115,16'h0016,16'h0113,-16'h00c0,-16'h00fc,-16'h00e3,16'h0019,16'h0071,-16'h0086,-16'h0070,16'h0004,16'h0022,16'h0000,-16'h003b,16'h0010,-16'h000c,-16'h000f,16'h000c,-16'h0001,16'h0010,-16'h0027,-16'h0029,16'h0018,16'h0003,-16'h0021,16'h0023,-16'h0004,16'h0074,-16'h001d,16'h0036,-16'h0022,-16'h0066,-16'h002b,16'h0003,-16'h0016,16'h000d,16'h0028,-16'h0036,16'h001c,-16'h0011,-16'h0017,-16'h0043,16'h003c,16'h0000,-16'h0018,-16'h000e,16'h0024,16'h0033,16'h0054,-16'h0058,16'h0032,16'h0030,16'h0032,-16'h0007,-16'h0024,-16'h0035,16'h003a,16'h0050,16'h002a,16'h0076,16'h0015,16'h000b,16'h0025,16'h000b,16'h005c,16'h000c,-16'h001c,-16'h0035,-16'h0063,16'h0016,-16'h000d,16'h0058,16'h0042,-16'h0060,-16'h0006,16'h0056,-16'h001d,16'h0027,-16'h004d,-16'h0031,-16'h0020,16'h0053,16'h002d,16'h005b,-16'h001d,16'h0022,16'h0093,-16'h0004,-16'h0019,16'h0007,-16'h004c,-16'h000b,-16'h0024,16'h0031,-16'h003c,-16'h000d,-16'h003d,16'h0008,16'h0032,-16'h0051,16'h0048,-16'h0070,-16'h004c,-16'h0013,-16'h0035,16'h000c,16'h010a,16'h0080,16'h0034,-16'h0038,16'h004d,-16'h0011,16'h0083,16'h0002,16'h003d,16'h0037,16'h0049,-16'h000b,16'h0007,16'h000d,16'h0015,-16'h0035,16'h0034,16'h000b,16'h0058,-16'h0056,16'h0002,-16'h0082,16'h0009,16'h003a,16'h0007,-16'h0078,-16'h0016,16'h001c,16'h000d,16'h002d,-16'h0048,16'h0003,16'h0076,16'h0094,-16'h003a,16'h0010,-16'h0029,-16'h0005,-16'h000f,16'h0004,-16'h0021,16'h008d,-16'h0022,16'h0011,16'h0081,16'h0062,16'h003e,-16'h0060,16'h0066,-16'h0011,-16'h0003,16'h0003,16'h0010,-16'h0005,-16'h003c,-16'h001b,16'h002b,-16'h0014,16'h0040,-16'h008e,16'h0024,16'h0002,-16'h002f,-16'h0075,16'h0185,16'h009b,16'h004b,16'h000a,16'h0049,-16'h0030,16'h00ae,-16'h0057,16'h003b,16'h0026,16'h0008,16'h0067,-16'h006a,16'h0080,16'h0005,16'h001e,-16'h0005,16'h009c,-16'h002a,-16'h004f,-16'h0002,-16'h001a,-16'h004e,16'h00a1,-16'h0020,-16'h004c,-16'h0092,-16'h0012,-16'h0057,16'h0051,-16'h000c,-16'h0041,-16'h0048,16'h00db,-16'h0029,16'h000d,-16'h0061,-16'h0019,16'h0067,-16'h0001,-16'h006f,16'h00f1,-16'h00a3,-16'h000a,16'h0081,16'h003d,-16'h002b,-16'h002f,-16'h000e,16'h0074,-16'h003a,-16'h0053,16'h0001,-16'h004b,-16'h0018,-16'h003a,16'h00cd,16'h000d,16'h0098,-16'h00b5,-16'h0043,-16'h001d,-16'h00a4,16'h0028,16'h0199,16'h008f,-16'h000b,-16'h005c,16'h001c,16'h0001,16'h00af,16'h0024,16'h0008,16'h003e,-16'h005e,16'h0033,-16'h00a2,16'h00ac,16'h0068,16'h006d,-16'h0035,16'h0077,16'h004d,-16'h00c5,16'h000b,-16'h004a,-16'h0093,16'h0081,-16'h0028,-16'h0041,-16'h0062,-16'h0050,-16'h00e0,-16'h0034,16'h0007,-16'h003d,-16'h001b,16'h00ff,-16'h001d,16'h0014,16'h0023,16'h003d,16'h00ab,-16'h0093,-16'h0066,16'h0103,-16'h00a7,-16'h00c9,16'h00a8,-16'h001c,-16'h0077,16'h00a5,16'h000c,16'h00bc,-16'h0043,-16'h0058,-16'h0070,-16'h004f,16'h0014,-16'h0057,16'h018e,16'h0020,16'h0102,-16'h0069,-16'h0015,-16'h000e,-16'h00c3,16'h0070,16'h018e,16'h0112,16'h005c,16'h0002,16'h0052,16'h0007,16'h00c4,16'h004a,16'h0057,16'h000f,-16'h004f,16'h009d,-16'h009f,16'h00ad,16'h0028,16'h0063,-16'h0004,16'h007b,-16'h007e,-16'h00e6,16'h0072,16'h002a,-16'h0074,-16'h002f,-16'h00ef,-16'h0013,-16'h0118,-16'h0095,-16'h00d4,16'h006f,16'h0019,-16'h008f,-16'h00c1,16'h0161,16'h0005,16'h0022,-16'h00a0,16'h000f,16'h003e,-16'h00b8,-16'h00ed,16'h0110,-16'h012e,-16'h0038,16'h013c,16'h0055,-16'h00d3,16'h00fd,16'h000a,16'h007c,-16'h00c9,-16'h0098,-16'h0051,-16'h00bc,-16'h0048,-16'h000d,16'h0118,-16'h001b,16'h0126,-16'h0091,16'h001b,-16'h0024,-16'h0183,16'h002c,16'h0142,16'h010a,-16'h0004,16'h0065,16'h0063,16'h008b,16'h015e,16'h0001,-16'h0039,16'h0052,-16'h008a,16'h001d,-16'h0107,16'h00fc,-16'h0097,16'h00b6,-16'h006d,16'h0054,-16'h0022,-16'h008d,16'h0036,-16'h0005,-16'h0129,-16'h0013,-16'h013b,16'h001f,-16'h010a,-16'h0078,-16'h0068,16'h0114,-16'h0015,-16'h0057,-16'h003b,16'h0179,16'h001b,16'h0018,-16'h0047,16'h0081,16'h0051,-16'h00e3,-16'h009f,16'h0061,-16'h0163,-16'h0035,16'h00c7,16'h0059,-16'h0143,16'h0158,-16'h0003,16'h0060,-16'h00fb,-16'h004e,-16'h006f,-16'h005c,-16'h00ca,-16'h0066,16'h0143,-16'h0018,16'h0160,-16'h0020,-16'h0089,16'h004f,-16'h01ba,-16'h001c,16'h010e,16'h010b,-16'h005e,16'h0024,-16'h0018,16'h00d9,16'h0102,16'h0032,-16'h007b,16'h00be,16'h005b,16'h003e,-16'h0105,16'h0023,-16'h0123,16'h0134,-16'h007f,-16'h0009,-16'h00d1,-16'h00e7,16'h0026,-16'h001b,-16'h00f4,-16'h0089,-16'h01c3,16'h00ee,-16'h00cf,-16'h00ac,-16'h00ff,16'h01b1,16'h0012,-16'h00b4,-16'h00be,16'h0153,16'h0069,-16'h000c,-16'h0077,16'h0099,16'h00ba,-16'h007b,-16'h008d,16'h0058,-16'h0130,16'h0051,16'h0134,16'h00fd,-16'h01ba,16'h00e3,-16'h000d,16'h00cf,-16'h018a,-16'h006a,-16'h0035,-16'h00cd,-16'h007b,16'h0002,16'h014d,-16'h0064,16'h0125,-16'h003f,-16'h00f0,-16'h0021,-16'h0144,-16'h000e,16'h0034,16'h014c,-16'h0018,16'h0018,-16'h0048,16'h0105,16'h0041,16'h0045,-16'h007d,16'h0114,16'h009c,16'h0015,-16'h005c,-16'h0015,-16'h00ce,16'h0147,16'h001d,16'h0002,-16'h00df,-16'h0180,16'h007a,-16'h0022,-16'h00cc,-16'h0061,-16'h0224,16'h0146,-16'h0171,-16'h00cf,-16'h00d8,16'h01dd,16'h0084,-16'h0084,16'h0009,16'h0121,16'h0026,-16'h00a2,-16'h007d,16'h0056,16'h0092,-16'h0085,-16'h0012,16'h001c,-16'h014d,16'h0102,16'h00d4,16'h0159,-16'h0197,16'h0008,-16'h0045,16'h0090,-16'h0249,16'h0085,16'h0011,-16'h007a,-16'h005c,16'h003b,16'h0205,-16'h006b,-16'h004d,-16'h000c,-16'h00ef,16'h003f,-16'h00ea,-16'h0022,-16'h0027,16'h0084,-16'h000b,-16'h0052,16'h0039,16'h012c,-16'h0011,-16'h00c0,-16'h0089,16'h00b7,16'h00aa,-16'h0073,16'h0043,-16'h0069,-16'h00cc,16'h01b1,-16'h0025,-16'h005d,-16'h00c4,-16'h015b,16'h010b,16'h0022,-16'h0108,-16'h00ac,-16'h01dd,16'h01d5,-16'h016c,-16'h0110,-16'h0050,16'h01a9,-16'h0006,-16'h0026,16'h0001,16'h016b,-16'h0073,-16'h0069,-16'h00ab,16'h0060,16'h007f,-16'h0092,16'h0037,16'h003c,-16'h00dd,16'h0139,16'h0075,16'h0160,-16'h0122,-16'h003d,16'h0014,16'h005b,-16'h0200,16'h001e,16'h00d6,16'h000a,-16'h002c,-16'h0003,16'h019b,-16'h002a,-16'h017c,16'h005e,-16'h0079,16'h0036,16'h006e,-16'h000a,16'h0007,-16'h0081,-16'h0084,16'h0000,16'h00cf,16'h005b,-16'h000f,-16'h013f,-16'h00b8,16'h00b0,16'h008e,-16'h000f,16'h0114,-16'h0087,-16'h010b,16'h0175,16'h0011,-16'h0082,-16'h00cb,-16'h00c9,16'h00d1,16'h00e2,-16'h00f9,-16'h0113,-16'h01f0,16'h0192,-16'h00be,-16'h0139,-16'h0007,16'h01af,-16'h002b,-16'h0061,-16'h004a,16'h0114,-16'h00bc,-16'h008f,-16'h006c,16'h0052,16'h00dc,-16'h0061,-16'h0016,16'h0077,-16'h00d0,16'h0128,16'h0008,16'h01b5,-16'h0140,-16'h00b7,-16'h00b9,-16'h001f,-16'h0074,16'h008c,16'h00e3,16'h0046,-16'h0017,16'h0041,16'h0162,-16'h001f,-16'h0215,16'h004d,-16'h0032,-16'h000e,16'h01ff,-16'h0071,-16'h0056,-16'h00d5,-16'h001e,-16'h0046,16'h00d3,-16'h0086,16'h0069,-16'h00e3,-16'h0055,16'h0061,16'h0056,16'h0056,16'h013d,-16'h005e,-16'h00a7,16'h001f,-16'h0074,-16'h00ae,-16'h00e3,-16'h009e,16'h00ab,16'h0087,-16'h008d,-16'h0135,-16'h0233,16'h0161,-16'h00e3,-16'h0106,16'h000c,16'h0106,-16'h00ed,-16'h0027,-16'h001f,16'h012f,-16'h0064,-16'h0065,-16'h0038,-16'h0031,16'h008c,-16'h0048,-16'h00a6,16'h0067,-16'h00b6,16'h0136,16'h000c,16'h0185,-16'h0189,16'h0019,-16'h00d1,-16'h0006,16'h011d,16'h007f,16'h00ef,16'h0023,-16'h0042,16'h0074,16'h00fd,-16'h0048,-16'h014e,-16'h00aa,16'h0014,16'h0049,16'h027b,16'h000c,-16'h00d0,-16'h016f,16'h0104,-16'h008c,16'h00f3,-16'h00ad,16'h001b,16'h0021,-16'h00a0,16'h008e,16'h0078,16'h0014,16'h020f,16'h0014,-16'h00af,16'h0029,-16'h000a,-16'h00a0,-16'h00dc,-16'h010b,16'h00e9,16'h0094,-16'h00ff,-16'h010b,-16'h0153,16'h00bf,-16'h0044,-16'h010d,-16'h0074,16'h0168,-16'h01d7,-16'h0044,16'h001b,16'h011b,-16'h004d,-16'h0054,-16'h0024,16'h003f,16'h00d3,16'h0029,-16'h0079,16'h0059,-16'h00d0,16'h0027,-16'h0168,16'h00fd,-16'h01c4,16'h0081,16'h0000,16'h0019,16'h016c,16'h005e,-16'h000b,-16'h0011,-16'h0024,16'h0129,16'h0089,-16'h0038,-16'h001c,-16'h0176,-16'h0001,-16'h0038,16'h01fe,16'h0076,-16'h0131,-16'h00f4,16'h009a,-16'h00df,16'h00cd,-16'h006a,16'h001e,16'h0065,-16'h00f1,16'h0043,16'h00c0,-16'h0037,16'h0215,-16'h0083,-16'h0059,16'h0014,-16'h0047,-16'h0064,-16'h01a4,-16'h00d6,16'h00ab,16'h00a9,-16'h0082,-16'h00be,-16'h0057,16'h0057,-16'h002a,-16'h0154,-16'h007b,16'h01b8,-16'h0156,-16'h009a,-16'h0022,16'h00f0,16'h003c,-16'h0038,16'h00b2,-16'h0032,16'h00b4,16'h0065,-16'h00f1,16'h004b,-16'h000a,16'h0085,-16'h0154,16'h0037,-16'h01ee,16'h001c,-16'h0049,16'h002b,16'h01bc,-16'h0052,-16'h0075,-16'h00cc,16'h00c6,16'h00e2,16'h0014,-16'h0001,16'h00ea,-16'h0226,16'h0064,-16'h008d,16'h01cb,16'h0066,-16'h01af,-16'h0083,16'h01b3,-16'h00f3,16'h007a,-16'h000b,-16'h0050,16'h0082,-16'h010c,16'h009d,16'h0034,-16'h0033,16'h0240,-16'h0084,16'h0041,-16'h0150,-16'h0016,16'h0014,-16'h0111,-16'h01e0,16'h0120,16'h00c2,-16'h0048,-16'h00a6,16'h0032,-16'h009c,16'h0022,-16'h01db,-16'h00f3,16'h011a,-16'h0159,-16'h00d7,16'h0000,16'h0148,16'h0001,-16'h0023,16'h0098,16'h0037,16'h0053,16'h00ba,-16'h0086,-16'h0077,-16'h0077,16'h00ef,-16'h00f1,-16'h007b,-16'h0266,16'h00ea,-16'h004c,-16'h0096,16'h00e6,-16'h0060,-16'h0062,-16'h00d7,16'h008f,16'h00dd,-16'h00e7,16'h0075,16'h01f0,-16'h022b,16'h00a9,-16'h0082,16'h01dd,16'h00a9,-16'h0103,16'h0001,16'h019f,-16'h0171,-16'h001b,16'h0099,16'h0001,16'h0156,-16'h0040,16'h0088,16'h006f,-16'h0040,16'h025b,-16'h0077,16'h005a,-16'h01df,16'h001d,16'h0006,-16'h00f5,-16'h027d,16'h00fe,16'h00bc,-16'h0017,-16'h0133,16'h007c,-16'h001f,16'h006b,-16'h02a3,-16'h00a8,16'h0014,-16'h018b,-16'h0133,-16'h0024,16'h00c5,16'h003e,16'h0003,16'h008b,16'h0010,16'h000d,16'h0124,-16'h0040,-16'h005d,16'h0019,16'h00a4,-16'h010c,-16'h0056,-16'h0257,16'h013f,-16'h004b,-16'h00cd,16'h00f8,-16'h011b,-16'h0145,-16'h006e,16'h004c,16'h00da,-16'h010a,16'h00ac,16'h01b9,-16'h01aa,16'h0069,-16'h00a2,16'h0090,16'h00bb,-16'h00c2,16'h0153,16'h015a,-16'h00ad,16'h0025,16'h01d1,-16'h00ed,16'h0156,-16'h005d,16'h0079,16'h00d2,-16'h0014,16'h0267,-16'h00fd,16'h004e,-16'h0127,16'h0003,-16'h0036,-16'h010b,-16'h029a,16'h0148,16'h00e0,-16'h00a4,-16'h016b,16'h00de,16'h0081,-16'h001f,-16'h02af,-16'h0067,-16'h0083,-16'h010b,-16'h0109,16'h00b6,16'h0123,16'h0068,16'h00d6,16'h00f6,16'h0059,16'h0057,16'h0132,16'h0004,16'h0015,16'h0084,16'h0093,-16'h00c2,-16'h009b,-16'h01fd,16'h0162,16'h0070,-16'h0161,16'h00d8,-16'h017f,-16'h00d3,-16'h0100,16'h0030,16'h0028,-16'h0080,16'h00ec,16'h00c8,-16'h0197,16'h0039,-16'h001f,-16'h0068,16'h00a9,-16'h005b,16'h0139,16'h00f1,-16'h00fe,16'h0081,16'h01e1,-16'h00ee,16'h01ae,-16'h0069,16'h00c8,16'h0074,16'h00cc,16'h0222,-16'h0018,16'h00b2,-16'h00e1,16'h0061,-16'h0082,-16'h00b8,-16'h02b8,16'h019b,16'h00d5,-16'h00f9,-16'h0141,16'h009e,16'h01c6,16'h0029,-16'h039c,16'h0000,-16'h0089,-16'h0036,-16'h012c,-16'h0033,16'h00e1,16'h0082,16'h0135,16'h00cc,16'h003d,16'h0003,16'h0176,-16'h002d,-16'h002e,16'h0039,16'h0075,-16'h0035,-16'h005c,-16'h0215,16'h0112,-16'h005f,-16'h0163,16'h003a,-16'h0257,-16'h0108,-16'h00a9,16'h002e,-16'h000e,-16'h0130,16'h007d,16'h00c3,-16'h0223,16'h00b8,-16'h00af,-16'h014a,16'h0083,16'h000e,16'h0105,16'h0187,-16'h0099,16'h007e,16'h0152,-16'h0127,-16'h003b,16'h0066,16'h00ae,16'h00bc,16'h00d7,16'h01ad,-16'h0026,16'h002e,-16'h00d9,16'h0099,-16'h004c,16'h0014,-16'h0181,16'h01ac,16'h00c5,-16'h010d,-16'h01a9,16'h00b9,16'h016a,16'h00a8,-16'h03fc,-16'h0060,-16'h00d4,16'h0057,-16'h0075,-16'h00f8,16'h0059,-16'h008c,16'h01d6,16'h00c3,16'h00f4,16'h0089,16'h0119,16'h000d,-16'h00a0,-16'h0073,16'h0069,-16'h0082,16'h00a8,-16'h01f5,16'h0167,-16'h00bf,-16'h0250,16'h0138,-16'h0233,-16'h01cb,-16'h00c1,16'h0007,-16'h00e5,-16'h012e,16'h00cd,16'h00b1,-16'h00ec,16'h005b,-16'h005b,-16'h0091,16'h007a,16'h0036,16'h009c,16'h00d7,16'h001b,16'h0105,16'h003d,-16'h0125,-16'h00ff,16'h00ef,16'h012f,16'h008f,16'h01fb,16'h013e,-16'h0010,-16'h0021,-16'h0158,16'h0043,-16'h000f,-16'h001f,-16'h011d,16'h018b,16'h003e,-16'h015b,-16'h0166,16'h0079,16'h0208,16'h0081,-16'h042e,-16'h00a5,-16'h015c,-16'h0036,-16'h0062,-16'h00e3,16'h00a6,-16'h011e,16'h01a2,16'h00e4,16'h007b,16'h002f,16'h009c,16'h0001,-16'h008f,16'h001a,-16'h00b7,-16'h0054,16'h00ef,-16'h023f,16'h01a6,-16'h006e,-16'h0258,16'h0144,-16'h0281,-16'h018c,-16'h0103,16'h00b2,-16'h00ff,-16'h00b2,16'h0065,16'h0030,-16'h00be,-16'h007d,-16'h008d,-16'h0034,16'h002e,16'h006c,16'h0015,16'h00f6,16'h009f,16'h018d,16'h0027,16'h0057,-16'h0185,16'h008a,16'h01e0,16'h0061,16'h01e5,16'h00f8,16'h0000,16'h0036,-16'h00e0,16'h005f,-16'h0086,-16'h007f,-16'h00a4,16'h0154,16'h0053,-16'h0118,-16'h0155,16'h002d,16'h0275,16'h00ec,-16'h03f7,-16'h00f9,-16'h01a5,-16'h0071,16'h00b7,-16'h00d3,16'h0026,-16'h0237,16'h019f,16'h013a,16'h0051,16'h0019,16'h000d,-16'h0037,-16'h008b,-16'h0062,-16'h00d7,16'h000d,16'h0117,-16'h0212,16'h019e,16'h0002,-16'h0204,16'h00a5,-16'h028d,-16'h0135,-16'h00ff,16'h0178,-16'h0086,-16'h0130,16'h009b,-16'h0029,-16'h00bc,-16'h02d7,16'h003f,16'h0016,16'h0028,-16'h006d,16'h000e,16'h00be,16'h014b,16'h0210,-16'h0024,16'h0049,-16'h0125,16'h01dc,16'h01d6,-16'h0018,16'h01f8,16'h00e3,-16'h000f,16'h0047,-16'h00ff,16'h002e,-16'h0088,-16'h00f5,-16'h0158,16'h0110,-16'h003b,-16'h0203,-16'h00f0,16'h005a,16'h01e1,16'h004f,-16'h03f4,-16'h00a5,-16'h02d0,-16'h0079,16'h0085,-16'h0002,-16'h002a,-16'h013e,16'h0161,16'h00d6,16'h0006,16'h0065,-16'h005b,-16'h0033,-16'h00bc,-16'h00bc,-16'h0172,16'h00b3,16'h0161,-16'h01fe,16'h008b,16'h0052,-16'h01f7,16'h0036,-16'h026c,-16'h00d5,-16'h012c,16'h0116,-16'h00a0,-16'h01c1,16'h00e1,-16'h0030,-16'h00fa,-16'h03df,16'h001c,16'h0069,16'h007a,-16'h0069,-16'h002f,16'h00f1,16'h01c3,16'h023b,-16'h0035,16'h00a5,-16'h0090,16'h01f3,16'h01e4,-16'h00e3,16'h01d5,16'h0068,-16'h0027,16'h00cd,-16'h0129,16'h0088,16'h000b,-16'h008e,-16'h010b,16'h013c,-16'h007d,-16'h01ed,-16'h0077,-16'h0004,16'h008d,16'h0043,-16'h03ae,-16'h0051,-16'h032c,16'h0013,16'h0096,16'h00d6,-16'h0075,-16'h00d0,16'h0090,16'h00cf,16'h0035,16'h0012,-16'h00d6,16'h0033,-16'h011a,-16'h00a6,-16'h00be,16'h00c1,16'h00f3,-16'h0276,16'h007b,16'h007e,-16'h0267,-16'h015b,-16'h0271,-16'h0030,-16'h0168,16'h011f,-16'h000c,-16'h023a,16'h0121,16'h0007,-16'h0141,-16'h0328,16'h0052,16'h00d9,16'h0041,-16'h00a3,16'h003b,16'h0125,16'h01fc,16'h0261,-16'h0040,16'h0105,16'h00bc,16'h01e7,16'h02dd,-16'h00d0,16'h0182,-16'h0017,-16'h002e,16'h0075,-16'h00e2,16'h0081,16'h003b,-16'h006f,-16'h00b2,16'h011e,16'h0001,-16'h0230,-16'h005a,-16'h000c,-16'h000f,-16'h0094,-16'h0354,16'h0013,-16'h02ce,16'h0079,16'h0157,16'h0065,-16'h0105,-16'h0013,16'h0052,16'h0081,16'h0016,16'h0096,-16'h00bc,16'h0076,-16'h00ec,-16'h0021,-16'h004e,16'h0127,16'h00d2,-16'h0242,16'h00f7,16'h0033,-16'h0189,-16'h00c9,-16'h0207,16'h0080,-16'h00ff,16'h0143,16'h001f,-16'h01e8,16'h017f,-16'h008e,-16'h016f,-16'h0164,-16'h003d,16'h00d7,-16'h00fc,-16'h0037,-16'h006d,16'h0118,16'h0196,16'h02a1,16'h0025,16'h0165,16'h0148,16'h0129,16'h02f6,-16'h0171,16'h0157,16'h001f,-16'h0021,16'h0054,-16'h0099,16'h001c,16'h008e,-16'h008f,16'h00f9,16'h015e,-16'h00a3,-16'h018a,-16'h0050,16'h003d,-16'h009c,-16'h010f,-16'h026f,16'h005b,-16'h01d5,16'h00b3,16'h00cf,16'h00cd,-16'h0181,-16'h0053,16'h0062,16'h0078,16'h0091,16'h00ce,-16'h0092,16'h0140,-16'h00e8,-16'h005b,-16'h0052,16'h01ca,16'h00a6,-16'h01da,16'h0081,16'h003a,-16'h00be,-16'h009a,-16'h01c8,16'h005c,-16'h007e,16'h00ec,16'h0050,-16'h018a,16'h0179,-16'h0107,-16'h010b,-16'h00ff,16'h0004,-16'h0006,-16'h01dc,-16'h003f,-16'h00b4,16'h0108,16'h01a4,16'h0162,16'h001c,16'h00b4,16'h0080,16'h0131,16'h02d9,-16'h0226,16'h0121,16'h0036,-16'h0070,16'h0033,-16'h00c4,16'h0041,16'h00e3,-16'h006a,16'h0196,16'h00c8,-16'h00a1,-16'h0152,-16'h005a,16'h0089,-16'h00f5,-16'h0172,-16'h029a,16'h0015,-16'h00d1,16'h0090,16'h008f,16'h00a6,-16'h019d,-16'h0045,-16'h0013,16'h001e,16'h00af,16'h00ab,-16'h009b,16'h00ca,-16'h0059,-16'h0019,-16'h0057,16'h0274,16'h00c8,-16'h021a,16'h007c,16'h005d,-16'h0088,16'h0041,-16'h0135,16'h0088,-16'h0061,16'h00f0,16'h00dc,-16'h012c,16'h00ed,-16'h0129,-16'h0084,-16'h0026,16'h0013,16'h0062,-16'h0171,-16'h0031,-16'h011c,16'h007b,16'h0078,16'h0148,16'h0094,16'h005a,16'h00db,16'h0039,16'h0222,-16'h0191,16'h0106,-16'h000c,-16'h0044,-16'h0048,-16'h003e,16'h0028,16'h00b9,-16'h00c5,16'h01cb,16'h0060,-16'h00b1,-16'h011b,-16'h000b,16'h0171,-16'h003e,-16'h012e,-16'h01e3,-16'h003a,-16'h005e,16'h00b2,16'h00e1,16'h0082,-16'h00ce,16'h0029,16'h0000,16'h003b,16'h006d,16'h0083,-16'h0025,16'h0161,-16'h003c,-16'h0032,-16'h00bb,16'h0240,16'h0002,-16'h01fc,16'h0075,-16'h0002,-16'h002e,16'h005c,-16'h00e0,16'h0088,16'h002e,16'h00a2,16'h00b0,-16'h0088,16'h00d4,-16'h00c0,-16'h0022,-16'h0013,16'h004d,-16'h0009,-16'h014f,-16'h0030,-16'h00be,-16'h000a,16'h004a,16'h0032,16'h0067,-16'h0006,16'h0098,-16'h0081,16'h01e6,-16'h015b,16'h0166,16'h0004,16'h000b,-16'h0017,-16'h000a,16'h007f,-16'h0062,-16'h0041,16'h01c4,16'h003e,-16'h0016,-16'h0072,16'h0013,16'h01e7,-16'h0069,-16'h010d,-16'h015d,-16'h0019,-16'h0056,-16'h0004,16'h0060,16'h0039,-16'h0076,16'h0065,16'h0040,16'h008c,16'h0033,16'h0010,16'h003c,16'h0160,16'h001d,16'h0044,-16'h001e,16'h01ae,16'h008a,-16'h017b,-16'h0033,-16'h001f,-16'h0017,16'h0047,-16'h0010,16'h0098,16'h0010,16'h002e,16'h005f,16'h000b,16'h0003,-16'h00b9,-16'h0058,16'h000d,16'h007b,-16'h005c,-16'h00bb,16'h003f,-16'h005b,-16'h0042,-16'h0039,16'h0055,16'h0072,-16'h0001,-16'h0023,-16'h008f,16'h017e,-16'h00a9,16'h0161,-16'h0017,-16'h000d,-16'h0072,-16'h0009,16'h004d,16'h0025,-16'h0099,16'h00f9,16'h005a,-16'h001c,-16'h0062,16'h000a,16'h0146,-16'h005d,-16'h00af,-16'h0118,16'h0063,16'h0034,-16'h0028,16'h002d};
    localparam [1023:0] bias_0 = {16'h01d3,-16'h0350,-16'h0066,-16'h00e9,-16'h00f8,16'h0254,16'h0018,-16'h028b,-16'h0724,-16'h04f9,16'h013f,16'h0326,-16'h0369,16'h0028,-16'h0068,16'h01ed,16'h0340,-16'h0519,16'h0451,-16'h005e,16'h0520,-16'h07a1,-16'h0187,-16'h004d,16'h00a9,-16'h02c3,16'h0075,16'h0002,16'h00ba,-16'h00ba,16'h043c,16'h0033,-16'h02fd,16'h02ec,-16'h00bb,16'h038e,16'h01d6,16'h0304,-16'h062a,16'h01b2,16'h0176,-16'h03a6,-16'h01ea,-16'h0401,16'h006e,-16'h00a3,-16'h022d,16'h0182,-16'h044a,16'h0261,-16'h00df,-16'h03f1,-16'h0701,16'h01c7,16'h01bd,-16'h03bd,-16'h03aa,-16'h01bd,-16'h0593,-16'h028a,-16'h05de,-16'h0418,16'h00fc,-16'h0124};

    localparam SWAIT = 3'd0;
    localparam SDOT = 3'd1;
    localparam SRELU = 3'd2;
    localparam SBIAS = 3'd3;
    localparam SFIN = 3'd4;
    reg [2:0] state, next_state;

    // row * WIDTH + col
    reg  [16 - 1:0] col, next_col;
    reg  [16*64 - 1:0] next_layer_0;
    reg  next_finish;

    always @(posedge clk ) begin
        if(rst) begin
            state <= SWAIT;
            col <= 0;
            layer_0 <= 0;
            finish <= 0;
        end else begin
            state <= next_state;
            col <= next_col;
            layer_0 <= next_layer_0;
            finish <= next_finish;
        end
    end
    // state
    always @(*) begin
        case (state)
            SWAIT: begin
                if(start) next_state = SDOT;
                else next_state = state;
            end
            SDOT: begin
                if(col == WIDTH - 1) next_state = SRELU;
                else next_state = state;
            end
            SRELU: next_state = SFIN;
            default: next_state = SWAIT;
        endcase
    end
    // row, col
    always @(*) begin
        case (state)
            SDOT: next_col = col + 16'b1;
            default: next_col = 16'b0;
        endcase
    end
    // finish
    always @(*) begin
        case (state)
            SBIAS: next_finish = 1'b1;
            default: next_finish = 1'b0;
        endcase
    end
    // layer_0
    always @(*) begin
        case (state)
            SWAIT: begin
                if(start) next_layer_0 = 0;
                else next_layer_0 = layer_0;
            end
            SDOT: begin
                next_layer_0[15-:16] = layer_0[15-:16] + layer_input[15-:16]*kernel_0[(0+col+1)*16-1-:16];
                next_layer_0[31-:16] = layer_0[31-:16] + layer_input[31-:16]*kernel_0[(64+col+1)*16-1-:16];
                next_layer_0[47-:16] = layer_0[47-:16] + layer_input[47-:16]*kernel_0[(128+col+1)*16-1-:16];
                next_layer_0[63-:16] = layer_0[63-:16] + layer_input[63-:16]*kernel_0[(192+col+1)*16-1-:16];
                next_layer_0[79-:16] = layer_0[79-:16] + layer_input[79-:16]*kernel_0[(256+col+1)*16-1-:16];
                next_layer_0[95-:16] = layer_0[95-:16] + layer_input[95-:16]*kernel_0[(320+col+1)*16-1-:16];
                next_layer_0[111-:16] = layer_0[111-:16] + layer_input[111-:16]*kernel_0[(384+col+1)*16-1-:16];
                next_layer_0[127-:16] = layer_0[127-:16] + layer_input[127-:16]*kernel_0[(448+col+1)*16-1-:16];
                next_layer_0[143-:16] = layer_0[143-:16] + layer_input[143-:16]*kernel_0[(512+col+1)*16-1-:16];
                next_layer_0[159-:16] = layer_0[159-:16] + layer_input[159-:16]*kernel_0[(576+col+1)*16-1-:16];
                next_layer_0[175-:16] = layer_0[175-:16] + layer_input[175-:16]*kernel_0[(640+col+1)*16-1-:16];
                next_layer_0[191-:16] = layer_0[191-:16] + layer_input[191-:16]*kernel_0[(704+col+1)*16-1-:16];
                next_layer_0[207-:16] = layer_0[207-:16] + layer_input[207-:16]*kernel_0[(768+col+1)*16-1-:16];
                next_layer_0[223-:16] = layer_0[223-:16] + layer_input[223-:16]*kernel_0[(832+col+1)*16-1-:16];
                next_layer_0[239-:16] = layer_0[239-:16] + layer_input[239-:16]*kernel_0[(896+col+1)*16-1-:16];
                next_layer_0[255-:16] = layer_0[255-:16] + layer_input[255-:16]*kernel_0[(960+col+1)*16-1-:16];
                next_layer_0[271-:16] = layer_0[271-:16] + layer_input[271-:16]*kernel_0[(1024+col+1)*16-1-:16];
                next_layer_0[287-:16] = layer_0[287-:16] + layer_input[287-:16]*kernel_0[(1088+col+1)*16-1-:16];
                next_layer_0[303-:16] = layer_0[303-:16] + layer_input[303-:16]*kernel_0[(1152+col+1)*16-1-:16];
                next_layer_0[319-:16] = layer_0[319-:16] + layer_input[319-:16]*kernel_0[(1216+col+1)*16-1-:16];
                next_layer_0[335-:16] = layer_0[335-:16] + layer_input[335-:16]*kernel_0[(1280+col+1)*16-1-:16];
                next_layer_0[351-:16] = layer_0[351-:16] + layer_input[351-:16]*kernel_0[(1344+col+1)*16-1-:16];
                next_layer_0[367-:16] = layer_0[367-:16] + layer_input[367-:16]*kernel_0[(1408+col+1)*16-1-:16];
                next_layer_0[383-:16] = layer_0[383-:16] + layer_input[383-:16]*kernel_0[(1472+col+1)*16-1-:16];
                next_layer_0[399-:16] = layer_0[399-:16] + layer_input[399-:16]*kernel_0[(1536+col+1)*16-1-:16];
                next_layer_0[415-:16] = layer_0[415-:16] + layer_input[415-:16]*kernel_0[(1600+col+1)*16-1-:16];
                next_layer_0[431-:16] = layer_0[431-:16] + layer_input[431-:16]*kernel_0[(1664+col+1)*16-1-:16];
                next_layer_0[447-:16] = layer_0[447-:16] + layer_input[447-:16]*kernel_0[(1728+col+1)*16-1-:16];
                next_layer_0[463-:16] = layer_0[463-:16] + layer_input[463-:16]*kernel_0[(1792+col+1)*16-1-:16];
                next_layer_0[479-:16] = layer_0[479-:16] + layer_input[479-:16]*kernel_0[(1856+col+1)*16-1-:16];
                next_layer_0[495-:16] = layer_0[495-:16] + layer_input[495-:16]*kernel_0[(1920+col+1)*16-1-:16];
                next_layer_0[511-:16] = layer_0[511-:16] + layer_input[511-:16]*kernel_0[(1984+col+1)*16-1-:16];
                next_layer_0[527-:16] = layer_0[527-:16] + layer_input[527-:16]*kernel_0[(2048+col+1)*16-1-:16];
                next_layer_0[543-:16] = layer_0[543-:16] + layer_input[543-:16]*kernel_0[(2112+col+1)*16-1-:16];
                next_layer_0[559-:16] = layer_0[559-:16] + layer_input[559-:16]*kernel_0[(2176+col+1)*16-1-:16];
                next_layer_0[575-:16] = layer_0[575-:16] + layer_input[575-:16]*kernel_0[(2240+col+1)*16-1-:16];
                next_layer_0[591-:16] = layer_0[591-:16] + layer_input[591-:16]*kernel_0[(2304+col+1)*16-1-:16];
                next_layer_0[607-:16] = layer_0[607-:16] + layer_input[607-:16]*kernel_0[(2368+col+1)*16-1-:16];
                next_layer_0[623-:16] = layer_0[623-:16] + layer_input[623-:16]*kernel_0[(2432+col+1)*16-1-:16];
                next_layer_0[639-:16] = layer_0[639-:16] + layer_input[639-:16]*kernel_0[(2496+col+1)*16-1-:16];
                next_layer_0[655-:16] = layer_0[655-:16] + layer_input[655-:16]*kernel_0[(2560+col+1)*16-1-:16];
                next_layer_0[671-:16] = layer_0[671-:16] + layer_input[671-:16]*kernel_0[(2624+col+1)*16-1-:16];
                next_layer_0[687-:16] = layer_0[687-:16] + layer_input[687-:16]*kernel_0[(2688+col+1)*16-1-:16];
                next_layer_0[703-:16] = layer_0[703-:16] + layer_input[703-:16]*kernel_0[(2752+col+1)*16-1-:16];
                next_layer_0[719-:16] = layer_0[719-:16] + layer_input[719-:16]*kernel_0[(2816+col+1)*16-1-:16];
                next_layer_0[735-:16] = layer_0[735-:16] + layer_input[735-:16]*kernel_0[(2880+col+1)*16-1-:16];
                next_layer_0[751-:16] = layer_0[751-:16] + layer_input[751-:16]*kernel_0[(2944+col+1)*16-1-:16];
                next_layer_0[767-:16] = layer_0[767-:16] + layer_input[767-:16]*kernel_0[(3008+col+1)*16-1-:16];
                next_layer_0[783-:16] = layer_0[783-:16] + layer_input[783-:16]*kernel_0[(3072+col+1)*16-1-:16];
                next_layer_0[799-:16] = layer_0[799-:16] + layer_input[799-:16]*kernel_0[(3136+col+1)*16-1-:16];
                next_layer_0[815-:16] = layer_0[815-:16] + layer_input[815-:16]*kernel_0[(3200+col+1)*16-1-:16];
                next_layer_0[831-:16] = layer_0[831-:16] + layer_input[831-:16]*kernel_0[(3264+col+1)*16-1-:16];
                next_layer_0[847-:16] = layer_0[847-:16] + layer_input[847-:16]*kernel_0[(3328+col+1)*16-1-:16];
                next_layer_0[863-:16] = layer_0[863-:16] + layer_input[863-:16]*kernel_0[(3392+col+1)*16-1-:16];
                next_layer_0[879-:16] = layer_0[879-:16] + layer_input[879-:16]*kernel_0[(3456+col+1)*16-1-:16];
                next_layer_0[895-:16] = layer_0[895-:16] + layer_input[895-:16]*kernel_0[(3520+col+1)*16-1-:16];
                next_layer_0[911-:16] = layer_0[911-:16] + layer_input[911-:16]*kernel_0[(3584+col+1)*16-1-:16];
                next_layer_0[927-:16] = layer_0[927-:16] + layer_input[927-:16]*kernel_0[(3648+col+1)*16-1-:16];
                next_layer_0[943-:16] = layer_0[943-:16] + layer_input[943-:16]*kernel_0[(3712+col+1)*16-1-:16];
                next_layer_0[959-:16] = layer_0[959-:16] + layer_input[959-:16]*kernel_0[(3776+col+1)*16-1-:16];
                next_layer_0[975-:16] = layer_0[975-:16] + layer_input[975-:16]*kernel_0[(3840+col+1)*16-1-:16];
                next_layer_0[991-:16] = layer_0[991-:16] + layer_input[991-:16]*kernel_0[(3904+col+1)*16-1-:16];
                next_layer_0[1007-:16] = layer_0[1007-:16] + layer_input[1007-:16]*kernel_0[(3968+col+1)*16-1-:16];
                next_layer_0[1023-:16] = layer_0[1023-:16] + layer_input[1023-:16]*kernel_0[(4032+col+1)*16-1-:16];
                next_layer_0[1039-:16] = layer_0[1039-:16] + layer_input[1039-:16]*kernel_0[(4096+col+1)*16-1-:16];
                next_layer_0[1055-:16] = layer_0[1055-:16] + layer_input[1055-:16]*kernel_0[(4160+col+1)*16-1-:16];
                next_layer_0[1071-:16] = layer_0[1071-:16] + layer_input[1071-:16]*kernel_0[(4224+col+1)*16-1-:16];
                next_layer_0[1087-:16] = layer_0[1087-:16] + layer_input[1087-:16]*kernel_0[(4288+col+1)*16-1-:16];
                next_layer_0[1103-:16] = layer_0[1103-:16] + layer_input[1103-:16]*kernel_0[(4352+col+1)*16-1-:16];
                next_layer_0[1119-:16] = layer_0[1119-:16] + layer_input[1119-:16]*kernel_0[(4416+col+1)*16-1-:16];
                next_layer_0[1135-:16] = layer_0[1135-:16] + layer_input[1135-:16]*kernel_0[(4480+col+1)*16-1-:16];
                next_layer_0[1151-:16] = layer_0[1151-:16] + layer_input[1151-:16]*kernel_0[(4544+col+1)*16-1-:16];
                next_layer_0[1167-:16] = layer_0[1167-:16] + layer_input[1167-:16]*kernel_0[(4608+col+1)*16-1-:16];
                next_layer_0[1183-:16] = layer_0[1183-:16] + layer_input[1183-:16]*kernel_0[(4672+col+1)*16-1-:16];
                next_layer_0[1199-:16] = layer_0[1199-:16] + layer_input[1199-:16]*kernel_0[(4736+col+1)*16-1-:16];
                next_layer_0[1215-:16] = layer_0[1215-:16] + layer_input[1215-:16]*kernel_0[(4800+col+1)*16-1-:16];
                next_layer_0[1231-:16] = layer_0[1231-:16] + layer_input[1231-:16]*kernel_0[(4864+col+1)*16-1-:16];
                next_layer_0[1247-:16] = layer_0[1247-:16] + layer_input[1247-:16]*kernel_0[(4928+col+1)*16-1-:16];
                next_layer_0[1263-:16] = layer_0[1263-:16] + layer_input[1263-:16]*kernel_0[(4992+col+1)*16-1-:16];
                next_layer_0[1279-:16] = layer_0[1279-:16] + layer_input[1279-:16]*kernel_0[(5056+col+1)*16-1-:16];
                next_layer_0[1295-:16] = layer_0[1295-:16] + layer_input[1295-:16]*kernel_0[(5120+col+1)*16-1-:16];
                next_layer_0[1311-:16] = layer_0[1311-:16] + layer_input[1311-:16]*kernel_0[(5184+col+1)*16-1-:16];
                next_layer_0[1327-:16] = layer_0[1327-:16] + layer_input[1327-:16]*kernel_0[(5248+col+1)*16-1-:16];
                next_layer_0[1343-:16] = layer_0[1343-:16] + layer_input[1343-:16]*kernel_0[(5312+col+1)*16-1-:16];
                next_layer_0[1359-:16] = layer_0[1359-:16] + layer_input[1359-:16]*kernel_0[(5376+col+1)*16-1-:16];
                next_layer_0[1375-:16] = layer_0[1375-:16] + layer_input[1375-:16]*kernel_0[(5440+col+1)*16-1-:16];
                next_layer_0[1391-:16] = layer_0[1391-:16] + layer_input[1391-:16]*kernel_0[(5504+col+1)*16-1-:16];
                next_layer_0[1407-:16] = layer_0[1407-:16] + layer_input[1407-:16]*kernel_0[(5568+col+1)*16-1-:16];
                next_layer_0[1423-:16] = layer_0[1423-:16] + layer_input[1423-:16]*kernel_0[(5632+col+1)*16-1-:16];
                next_layer_0[1439-:16] = layer_0[1439-:16] + layer_input[1439-:16]*kernel_0[(5696+col+1)*16-1-:16];
                next_layer_0[1455-:16] = layer_0[1455-:16] + layer_input[1455-:16]*kernel_0[(5760+col+1)*16-1-:16];
                next_layer_0[1471-:16] = layer_0[1471-:16] + layer_input[1471-:16]*kernel_0[(5824+col+1)*16-1-:16];
                next_layer_0[1487-:16] = layer_0[1487-:16] + layer_input[1487-:16]*kernel_0[(5888+col+1)*16-1-:16];
                next_layer_0[1503-:16] = layer_0[1503-:16] + layer_input[1503-:16]*kernel_0[(5952+col+1)*16-1-:16];
                next_layer_0[1519-:16] = layer_0[1519-:16] + layer_input[1519-:16]*kernel_0[(6016+col+1)*16-1-:16];
                next_layer_0[1535-:16] = layer_0[1535-:16] + layer_input[1535-:16]*kernel_0[(6080+col+1)*16-1-:16];
                next_layer_0[1551-:16] = layer_0[1551-:16] + layer_input[1551-:16]*kernel_0[(6144+col+1)*16-1-:16];
                next_layer_0[1567-:16] = layer_0[1567-:16] + layer_input[1567-:16]*kernel_0[(6208+col+1)*16-1-:16];
                next_layer_0[1583-:16] = layer_0[1583-:16] + layer_input[1583-:16]*kernel_0[(6272+col+1)*16-1-:16];
                next_layer_0[1599-:16] = layer_0[1599-:16] + layer_input[1599-:16]*kernel_0[(6336+col+1)*16-1-:16];
                next_layer_0[1615-:16] = layer_0[1615-:16] + layer_input[1615-:16]*kernel_0[(6400+col+1)*16-1-:16];
                next_layer_0[1631-:16] = layer_0[1631-:16] + layer_input[1631-:16]*kernel_0[(6464+col+1)*16-1-:16];
                next_layer_0[1647-:16] = layer_0[1647-:16] + layer_input[1647-:16]*kernel_0[(6528+col+1)*16-1-:16];
                next_layer_0[1663-:16] = layer_0[1663-:16] + layer_input[1663-:16]*kernel_0[(6592+col+1)*16-1-:16];
                next_layer_0[1679-:16] = layer_0[1679-:16] + layer_input[1679-:16]*kernel_0[(6656+col+1)*16-1-:16];
                next_layer_0[1695-:16] = layer_0[1695-:16] + layer_input[1695-:16]*kernel_0[(6720+col+1)*16-1-:16];
                next_layer_0[1711-:16] = layer_0[1711-:16] + layer_input[1711-:16]*kernel_0[(6784+col+1)*16-1-:16];
                next_layer_0[1727-:16] = layer_0[1727-:16] + layer_input[1727-:16]*kernel_0[(6848+col+1)*16-1-:16];
                next_layer_0[1743-:16] = layer_0[1743-:16] + layer_input[1743-:16]*kernel_0[(6912+col+1)*16-1-:16];
                next_layer_0[1759-:16] = layer_0[1759-:16] + layer_input[1759-:16]*kernel_0[(6976+col+1)*16-1-:16];
                next_layer_0[1775-:16] = layer_0[1775-:16] + layer_input[1775-:16]*kernel_0[(7040+col+1)*16-1-:16];
                next_layer_0[1791-:16] = layer_0[1791-:16] + layer_input[1791-:16]*kernel_0[(7104+col+1)*16-1-:16];
                next_layer_0[1807-:16] = layer_0[1807-:16] + layer_input[1807-:16]*kernel_0[(7168+col+1)*16-1-:16];
                next_layer_0[1823-:16] = layer_0[1823-:16] + layer_input[1823-:16]*kernel_0[(7232+col+1)*16-1-:16];
                next_layer_0[1839-:16] = layer_0[1839-:16] + layer_input[1839-:16]*kernel_0[(7296+col+1)*16-1-:16];
                next_layer_0[1855-:16] = layer_0[1855-:16] + layer_input[1855-:16]*kernel_0[(7360+col+1)*16-1-:16];
                next_layer_0[1871-:16] = layer_0[1871-:16] + layer_input[1871-:16]*kernel_0[(7424+col+1)*16-1-:16];
                next_layer_0[1887-:16] = layer_0[1887-:16] + layer_input[1887-:16]*kernel_0[(7488+col+1)*16-1-:16];
                next_layer_0[1903-:16] = layer_0[1903-:16] + layer_input[1903-:16]*kernel_0[(7552+col+1)*16-1-:16];
                next_layer_0[1919-:16] = layer_0[1919-:16] + layer_input[1919-:16]*kernel_0[(7616+col+1)*16-1-:16];
                next_layer_0[1935-:16] = layer_0[1935-:16] + layer_input[1935-:16]*kernel_0[(7680+col+1)*16-1-:16];
                next_layer_0[1951-:16] = layer_0[1951-:16] + layer_input[1951-:16]*kernel_0[(7744+col+1)*16-1-:16];
                next_layer_0[1967-:16] = layer_0[1967-:16] + layer_input[1967-:16]*kernel_0[(7808+col+1)*16-1-:16];
                next_layer_0[1983-:16] = layer_0[1983-:16] + layer_input[1983-:16]*kernel_0[(7872+col+1)*16-1-:16];
                next_layer_0[1999-:16] = layer_0[1999-:16] + layer_input[1999-:16]*kernel_0[(7936+col+1)*16-1-:16];
                next_layer_0[2015-:16] = layer_0[2015-:16] + layer_input[2015-:16]*kernel_0[(8000+col+1)*16-1-:16];
                next_layer_0[2031-:16] = layer_0[2031-:16] + layer_input[2031-:16]*kernel_0[(8064+col+1)*16-1-:16];
                next_layer_0[2047-:16] = layer_0[2047-:16] + layer_input[2047-:16]*kernel_0[(8128+col+1)*16-1-:16];
                next_layer_0[2063-:16] = layer_0[2063-:16] + layer_input[2063-:16]*kernel_0[(8192+col+1)*16-1-:16];
                next_layer_0[2079-:16] = layer_0[2079-:16] + layer_input[2079-:16]*kernel_0[(8256+col+1)*16-1-:16];
                next_layer_0[2095-:16] = layer_0[2095-:16] + layer_input[2095-:16]*kernel_0[(8320+col+1)*16-1-:16];
                next_layer_0[2111-:16] = layer_0[2111-:16] + layer_input[2111-:16]*kernel_0[(8384+col+1)*16-1-:16];
                next_layer_0[2127-:16] = layer_0[2127-:16] + layer_input[2127-:16]*kernel_0[(8448+col+1)*16-1-:16];
                next_layer_0[2143-:16] = layer_0[2143-:16] + layer_input[2143-:16]*kernel_0[(8512+col+1)*16-1-:16];
                next_layer_0[2159-:16] = layer_0[2159-:16] + layer_input[2159-:16]*kernel_0[(8576+col+1)*16-1-:16];
                next_layer_0[2175-:16] = layer_0[2175-:16] + layer_input[2175-:16]*kernel_0[(8640+col+1)*16-1-:16];
                next_layer_0[2191-:16] = layer_0[2191-:16] + layer_input[2191-:16]*kernel_0[(8704+col+1)*16-1-:16];
                next_layer_0[2207-:16] = layer_0[2207-:16] + layer_input[2207-:16]*kernel_0[(8768+col+1)*16-1-:16];
                next_layer_0[2223-:16] = layer_0[2223-:16] + layer_input[2223-:16]*kernel_0[(8832+col+1)*16-1-:16];
                next_layer_0[2239-:16] = layer_0[2239-:16] + layer_input[2239-:16]*kernel_0[(8896+col+1)*16-1-:16];
                next_layer_0[2255-:16] = layer_0[2255-:16] + layer_input[2255-:16]*kernel_0[(8960+col+1)*16-1-:16];
                next_layer_0[2271-:16] = layer_0[2271-:16] + layer_input[2271-:16]*kernel_0[(9024+col+1)*16-1-:16];
                next_layer_0[2287-:16] = layer_0[2287-:16] + layer_input[2287-:16]*kernel_0[(9088+col+1)*16-1-:16];
                next_layer_0[2303-:16] = layer_0[2303-:16] + layer_input[2303-:16]*kernel_0[(9152+col+1)*16-1-:16];
                next_layer_0[2319-:16] = layer_0[2319-:16] + layer_input[2319-:16]*kernel_0[(9216+col+1)*16-1-:16];
                next_layer_0[2335-:16] = layer_0[2335-:16] + layer_input[2335-:16]*kernel_0[(9280+col+1)*16-1-:16];
                next_layer_0[2351-:16] = layer_0[2351-:16] + layer_input[2351-:16]*kernel_0[(9344+col+1)*16-1-:16];
                next_layer_0[2367-:16] = layer_0[2367-:16] + layer_input[2367-:16]*kernel_0[(9408+col+1)*16-1-:16];
                next_layer_0[2383-:16] = layer_0[2383-:16] + layer_input[2383-:16]*kernel_0[(9472+col+1)*16-1-:16];
                next_layer_0[2399-:16] = layer_0[2399-:16] + layer_input[2399-:16]*kernel_0[(9536+col+1)*16-1-:16];
                next_layer_0[2415-:16] = layer_0[2415-:16] + layer_input[2415-:16]*kernel_0[(9600+col+1)*16-1-:16];
                next_layer_0[2431-:16] = layer_0[2431-:16] + layer_input[2431-:16]*kernel_0[(9664+col+1)*16-1-:16];
                next_layer_0[2447-:16] = layer_0[2447-:16] + layer_input[2447-:16]*kernel_0[(9728+col+1)*16-1-:16];
                next_layer_0[2463-:16] = layer_0[2463-:16] + layer_input[2463-:16]*kernel_0[(9792+col+1)*16-1-:16];
                next_layer_0[2479-:16] = layer_0[2479-:16] + layer_input[2479-:16]*kernel_0[(9856+col+1)*16-1-:16];
                next_layer_0[2495-:16] = layer_0[2495-:16] + layer_input[2495-:16]*kernel_0[(9920+col+1)*16-1-:16];
                next_layer_0[2511-:16] = layer_0[2511-:16] + layer_input[2511-:16]*kernel_0[(9984+col+1)*16-1-:16];
                next_layer_0[2527-:16] = layer_0[2527-:16] + layer_input[2527-:16]*kernel_0[(10048+col+1)*16-1-:16];
                next_layer_0[2543-:16] = layer_0[2543-:16] + layer_input[2543-:16]*kernel_0[(10112+col+1)*16-1-:16];
                next_layer_0[2559-:16] = layer_0[2559-:16] + layer_input[2559-:16]*kernel_0[(10176+col+1)*16-1-:16];
                next_layer_0[2575-:16] = layer_0[2575-:16] + layer_input[2575-:16]*kernel_0[(10240+col+1)*16-1-:16];
                next_layer_0[2591-:16] = layer_0[2591-:16] + layer_input[2591-:16]*kernel_0[(10304+col+1)*16-1-:16];
                next_layer_0[2607-:16] = layer_0[2607-:16] + layer_input[2607-:16]*kernel_0[(10368+col+1)*16-1-:16];
                next_layer_0[2623-:16] = layer_0[2623-:16] + layer_input[2623-:16]*kernel_0[(10432+col+1)*16-1-:16];
                next_layer_0[2639-:16] = layer_0[2639-:16] + layer_input[2639-:16]*kernel_0[(10496+col+1)*16-1-:16];
                next_layer_0[2655-:16] = layer_0[2655-:16] + layer_input[2655-:16]*kernel_0[(10560+col+1)*16-1-:16];
                next_layer_0[2671-:16] = layer_0[2671-:16] + layer_input[2671-:16]*kernel_0[(10624+col+1)*16-1-:16];
                next_layer_0[2687-:16] = layer_0[2687-:16] + layer_input[2687-:16]*kernel_0[(10688+col+1)*16-1-:16];
                next_layer_0[2703-:16] = layer_0[2703-:16] + layer_input[2703-:16]*kernel_0[(10752+col+1)*16-1-:16];
                next_layer_0[2719-:16] = layer_0[2719-:16] + layer_input[2719-:16]*kernel_0[(10816+col+1)*16-1-:16];
                next_layer_0[2735-:16] = layer_0[2735-:16] + layer_input[2735-:16]*kernel_0[(10880+col+1)*16-1-:16];
                next_layer_0[2751-:16] = layer_0[2751-:16] + layer_input[2751-:16]*kernel_0[(10944+col+1)*16-1-:16];
                next_layer_0[2767-:16] = layer_0[2767-:16] + layer_input[2767-:16]*kernel_0[(11008+col+1)*16-1-:16];
                next_layer_0[2783-:16] = layer_0[2783-:16] + layer_input[2783-:16]*kernel_0[(11072+col+1)*16-1-:16];
                next_layer_0[2799-:16] = layer_0[2799-:16] + layer_input[2799-:16]*kernel_0[(11136+col+1)*16-1-:16];
                next_layer_0[2815-:16] = layer_0[2815-:16] + layer_input[2815-:16]*kernel_0[(11200+col+1)*16-1-:16];
                next_layer_0[2831-:16] = layer_0[2831-:16] + layer_input[2831-:16]*kernel_0[(11264+col+1)*16-1-:16];
                next_layer_0[2847-:16] = layer_0[2847-:16] + layer_input[2847-:16]*kernel_0[(11328+col+1)*16-1-:16];
                next_layer_0[2863-:16] = layer_0[2863-:16] + layer_input[2863-:16]*kernel_0[(11392+col+1)*16-1-:16];
                next_layer_0[2879-:16] = layer_0[2879-:16] + layer_input[2879-:16]*kernel_0[(11456+col+1)*16-1-:16];
                next_layer_0[2895-:16] = layer_0[2895-:16] + layer_input[2895-:16]*kernel_0[(11520+col+1)*16-1-:16];
                next_layer_0[2911-:16] = layer_0[2911-:16] + layer_input[2911-:16]*kernel_0[(11584+col+1)*16-1-:16];
                next_layer_0[2927-:16] = layer_0[2927-:16] + layer_input[2927-:16]*kernel_0[(11648+col+1)*16-1-:16];
                next_layer_0[2943-:16] = layer_0[2943-:16] + layer_input[2943-:16]*kernel_0[(11712+col+1)*16-1-:16];
                next_layer_0[2959-:16] = layer_0[2959-:16] + layer_input[2959-:16]*kernel_0[(11776+col+1)*16-1-:16];
                next_layer_0[2975-:16] = layer_0[2975-:16] + layer_input[2975-:16]*kernel_0[(11840+col+1)*16-1-:16];
                next_layer_0[2991-:16] = layer_0[2991-:16] + layer_input[2991-:16]*kernel_0[(11904+col+1)*16-1-:16];
                next_layer_0[3007-:16] = layer_0[3007-:16] + layer_input[3007-:16]*kernel_0[(11968+col+1)*16-1-:16];
                next_layer_0[3023-:16] = layer_0[3023-:16] + layer_input[3023-:16]*kernel_0[(12032+col+1)*16-1-:16];
                next_layer_0[3039-:16] = layer_0[3039-:16] + layer_input[3039-:16]*kernel_0[(12096+col+1)*16-1-:16];
                next_layer_0[3055-:16] = layer_0[3055-:16] + layer_input[3055-:16]*kernel_0[(12160+col+1)*16-1-:16];
                next_layer_0[3071-:16] = layer_0[3071-:16] + layer_input[3071-:16]*kernel_0[(12224+col+1)*16-1-:16];
                next_layer_0[3087-:16] = layer_0[3087-:16] + layer_input[3087-:16]*kernel_0[(12288+col+1)*16-1-:16];
                next_layer_0[3103-:16] = layer_0[3103-:16] + layer_input[3103-:16]*kernel_0[(12352+col+1)*16-1-:16];
                next_layer_0[3119-:16] = layer_0[3119-:16] + layer_input[3119-:16]*kernel_0[(12416+col+1)*16-1-:16];
                next_layer_0[3135-:16] = layer_0[3135-:16] + layer_input[3135-:16]*kernel_0[(12480+col+1)*16-1-:16];
                next_layer_0[3151-:16] = layer_0[3151-:16] + layer_input[3151-:16]*kernel_0[(12544+col+1)*16-1-:16];
                next_layer_0[3167-:16] = layer_0[3167-:16] + layer_input[3167-:16]*kernel_0[(12608+col+1)*16-1-:16];
                next_layer_0[3183-:16] = layer_0[3183-:16] + layer_input[3183-:16]*kernel_0[(12672+col+1)*16-1-:16];
                next_layer_0[3199-:16] = layer_0[3199-:16] + layer_input[3199-:16]*kernel_0[(12736+col+1)*16-1-:16];
                next_layer_0[3215-:16] = layer_0[3215-:16] + layer_input[3215-:16]*kernel_0[(12800+col+1)*16-1-:16];
                next_layer_0[3231-:16] = layer_0[3231-:16] + layer_input[3231-:16]*kernel_0[(12864+col+1)*16-1-:16];
                next_layer_0[3247-:16] = layer_0[3247-:16] + layer_input[3247-:16]*kernel_0[(12928+col+1)*16-1-:16];
                next_layer_0[3263-:16] = layer_0[3263-:16] + layer_input[3263-:16]*kernel_0[(12992+col+1)*16-1-:16];
                next_layer_0[3279-:16] = layer_0[3279-:16] + layer_input[3279-:16]*kernel_0[(13056+col+1)*16-1-:16];
                next_layer_0[3295-:16] = layer_0[3295-:16] + layer_input[3295-:16]*kernel_0[(13120+col+1)*16-1-:16];
                next_layer_0[3311-:16] = layer_0[3311-:16] + layer_input[3311-:16]*kernel_0[(13184+col+1)*16-1-:16];
                next_layer_0[3327-:16] = layer_0[3327-:16] + layer_input[3327-:16]*kernel_0[(13248+col+1)*16-1-:16];
                next_layer_0[3343-:16] = layer_0[3343-:16] + layer_input[3343-:16]*kernel_0[(13312+col+1)*16-1-:16];
                next_layer_0[3359-:16] = layer_0[3359-:16] + layer_input[3359-:16]*kernel_0[(13376+col+1)*16-1-:16];
                next_layer_0[3375-:16] = layer_0[3375-:16] + layer_input[3375-:16]*kernel_0[(13440+col+1)*16-1-:16];
                next_layer_0[3391-:16] = layer_0[3391-:16] + layer_input[3391-:16]*kernel_0[(13504+col+1)*16-1-:16];
                next_layer_0[3407-:16] = layer_0[3407-:16] + layer_input[3407-:16]*kernel_0[(13568+col+1)*16-1-:16];
                next_layer_0[3423-:16] = layer_0[3423-:16] + layer_input[3423-:16]*kernel_0[(13632+col+1)*16-1-:16];
                next_layer_0[3439-:16] = layer_0[3439-:16] + layer_input[3439-:16]*kernel_0[(13696+col+1)*16-1-:16];
                next_layer_0[3455-:16] = layer_0[3455-:16] + layer_input[3455-:16]*kernel_0[(13760+col+1)*16-1-:16];
                next_layer_0[3471-:16] = layer_0[3471-:16] + layer_input[3471-:16]*kernel_0[(13824+col+1)*16-1-:16];
                next_layer_0[3487-:16] = layer_0[3487-:16] + layer_input[3487-:16]*kernel_0[(13888+col+1)*16-1-:16];
                next_layer_0[3503-:16] = layer_0[3503-:16] + layer_input[3503-:16]*kernel_0[(13952+col+1)*16-1-:16];
                next_layer_0[3519-:16] = layer_0[3519-:16] + layer_input[3519-:16]*kernel_0[(14016+col+1)*16-1-:16];
                next_layer_0[3535-:16] = layer_0[3535-:16] + layer_input[3535-:16]*kernel_0[(14080+col+1)*16-1-:16];
                next_layer_0[3551-:16] = layer_0[3551-:16] + layer_input[3551-:16]*kernel_0[(14144+col+1)*16-1-:16];
                next_layer_0[3567-:16] = layer_0[3567-:16] + layer_input[3567-:16]*kernel_0[(14208+col+1)*16-1-:16];
                next_layer_0[3583-:16] = layer_0[3583-:16] + layer_input[3583-:16]*kernel_0[(14272+col+1)*16-1-:16];
                next_layer_0[3599-:16] = layer_0[3599-:16] + layer_input[3599-:16]*kernel_0[(14336+col+1)*16-1-:16];
                next_layer_0[3615-:16] = layer_0[3615-:16] + layer_input[3615-:16]*kernel_0[(14400+col+1)*16-1-:16];
                next_layer_0[3631-:16] = layer_0[3631-:16] + layer_input[3631-:16]*kernel_0[(14464+col+1)*16-1-:16];
                next_layer_0[3647-:16] = layer_0[3647-:16] + layer_input[3647-:16]*kernel_0[(14528+col+1)*16-1-:16];
                next_layer_0[3663-:16] = layer_0[3663-:16] + layer_input[3663-:16]*kernel_0[(14592+col+1)*16-1-:16];
                next_layer_0[3679-:16] = layer_0[3679-:16] + layer_input[3679-:16]*kernel_0[(14656+col+1)*16-1-:16];
                next_layer_0[3695-:16] = layer_0[3695-:16] + layer_input[3695-:16]*kernel_0[(14720+col+1)*16-1-:16];
                next_layer_0[3711-:16] = layer_0[3711-:16] + layer_input[3711-:16]*kernel_0[(14784+col+1)*16-1-:16];
                next_layer_0[3727-:16] = layer_0[3727-:16] + layer_input[3727-:16]*kernel_0[(14848+col+1)*16-1-:16];
                next_layer_0[3743-:16] = layer_0[3743-:16] + layer_input[3743-:16]*kernel_0[(14912+col+1)*16-1-:16];
                next_layer_0[3759-:16] = layer_0[3759-:16] + layer_input[3759-:16]*kernel_0[(14976+col+1)*16-1-:16];
                next_layer_0[3775-:16] = layer_0[3775-:16] + layer_input[3775-:16]*kernel_0[(15040+col+1)*16-1-:16];
                next_layer_0[3791-:16] = layer_0[3791-:16] + layer_input[3791-:16]*kernel_0[(15104+col+1)*16-1-:16];
                next_layer_0[3807-:16] = layer_0[3807-:16] + layer_input[3807-:16]*kernel_0[(15168+col+1)*16-1-:16];
                next_layer_0[3823-:16] = layer_0[3823-:16] + layer_input[3823-:16]*kernel_0[(15232+col+1)*16-1-:16];
                next_layer_0[3839-:16] = layer_0[3839-:16] + layer_input[3839-:16]*kernel_0[(15296+col+1)*16-1-:16];
                next_layer_0[3855-:16] = layer_0[3855-:16] + layer_input[3855-:16]*kernel_0[(15360+col+1)*16-1-:16];
                next_layer_0[3871-:16] = layer_0[3871-:16] + layer_input[3871-:16]*kernel_0[(15424+col+1)*16-1-:16];
                next_layer_0[3887-:16] = layer_0[3887-:16] + layer_input[3887-:16]*kernel_0[(15488+col+1)*16-1-:16];
                next_layer_0[3903-:16] = layer_0[3903-:16] + layer_input[3903-:16]*kernel_0[(15552+col+1)*16-1-:16];
                next_layer_0[3919-:16] = layer_0[3919-:16] + layer_input[3919-:16]*kernel_0[(15616+col+1)*16-1-:16];
                next_layer_0[3935-:16] = layer_0[3935-:16] + layer_input[3935-:16]*kernel_0[(15680+col+1)*16-1-:16];
                next_layer_0[3951-:16] = layer_0[3951-:16] + layer_input[3951-:16]*kernel_0[(15744+col+1)*16-1-:16];
                next_layer_0[3967-:16] = layer_0[3967-:16] + layer_input[3967-:16]*kernel_0[(15808+col+1)*16-1-:16];
                next_layer_0[3983-:16] = layer_0[3983-:16] + layer_input[3983-:16]*kernel_0[(15872+col+1)*16-1-:16];
                next_layer_0[3999-:16] = layer_0[3999-:16] + layer_input[3999-:16]*kernel_0[(15936+col+1)*16-1-:16];
                next_layer_0[4015-:16] = layer_0[4015-:16] + layer_input[4015-:16]*kernel_0[(16000+col+1)*16-1-:16];
                next_layer_0[4031-:16] = layer_0[4031-:16] + layer_input[4031-:16]*kernel_0[(16064+col+1)*16-1-:16];
                next_layer_0[4047-:16] = layer_0[4047-:16] + layer_input[4047-:16]*kernel_0[(16128+col+1)*16-1-:16];
                next_layer_0[4063-:16] = layer_0[4063-:16] + layer_input[4063-:16]*kernel_0[(16192+col+1)*16-1-:16];
                next_layer_0[4079-:16] = layer_0[4079-:16] + layer_input[4079-:16]*kernel_0[(16256+col+1)*16-1-:16];
                next_layer_0[4095-:16] = layer_0[4095-:16] + layer_input[4095-:16]*kernel_0[(16320+col+1)*16-1-:16];
                next_layer_0[4111-:16] = layer_0[4111-:16] + layer_input[4111-:16]*kernel_0[(16384+col+1)*16-1-:16];
                next_layer_0[4127-:16] = layer_0[4127-:16] + layer_input[4127-:16]*kernel_0[(16448+col+1)*16-1-:16];
                next_layer_0[4143-:16] = layer_0[4143-:16] + layer_input[4143-:16]*kernel_0[(16512+col+1)*16-1-:16];
                next_layer_0[4159-:16] = layer_0[4159-:16] + layer_input[4159-:16]*kernel_0[(16576+col+1)*16-1-:16];
                next_layer_0[4175-:16] = layer_0[4175-:16] + layer_input[4175-:16]*kernel_0[(16640+col+1)*16-1-:16];
                next_layer_0[4191-:16] = layer_0[4191-:16] + layer_input[4191-:16]*kernel_0[(16704+col+1)*16-1-:16];
                next_layer_0[4207-:16] = layer_0[4207-:16] + layer_input[4207-:16]*kernel_0[(16768+col+1)*16-1-:16];
                next_layer_0[4223-:16] = layer_0[4223-:16] + layer_input[4223-:16]*kernel_0[(16832+col+1)*16-1-:16];
                next_layer_0[4239-:16] = layer_0[4239-:16] + layer_input[4239-:16]*kernel_0[(16896+col+1)*16-1-:16];
                next_layer_0[4255-:16] = layer_0[4255-:16] + layer_input[4255-:16]*kernel_0[(16960+col+1)*16-1-:16];
                next_layer_0[4271-:16] = layer_0[4271-:16] + layer_input[4271-:16]*kernel_0[(17024+col+1)*16-1-:16];
                next_layer_0[4287-:16] = layer_0[4287-:16] + layer_input[4287-:16]*kernel_0[(17088+col+1)*16-1-:16];
                next_layer_0[4303-:16] = layer_0[4303-:16] + layer_input[4303-:16]*kernel_0[(17152+col+1)*16-1-:16];
                next_layer_0[4319-:16] = layer_0[4319-:16] + layer_input[4319-:16]*kernel_0[(17216+col+1)*16-1-:16];
                next_layer_0[4335-:16] = layer_0[4335-:16] + layer_input[4335-:16]*kernel_0[(17280+col+1)*16-1-:16];
                next_layer_0[4351-:16] = layer_0[4351-:16] + layer_input[4351-:16]*kernel_0[(17344+col+1)*16-1-:16];
                next_layer_0[4367-:16] = layer_0[4367-:16] + layer_input[4367-:16]*kernel_0[(17408+col+1)*16-1-:16];
                next_layer_0[4383-:16] = layer_0[4383-:16] + layer_input[4383-:16]*kernel_0[(17472+col+1)*16-1-:16];
                next_layer_0[4399-:16] = layer_0[4399-:16] + layer_input[4399-:16]*kernel_0[(17536+col+1)*16-1-:16];
                next_layer_0[4415-:16] = layer_0[4415-:16] + layer_input[4415-:16]*kernel_0[(17600+col+1)*16-1-:16];
                next_layer_0[4431-:16] = layer_0[4431-:16] + layer_input[4431-:16]*kernel_0[(17664+col+1)*16-1-:16];
                next_layer_0[4447-:16] = layer_0[4447-:16] + layer_input[4447-:16]*kernel_0[(17728+col+1)*16-1-:16];
                next_layer_0[4463-:16] = layer_0[4463-:16] + layer_input[4463-:16]*kernel_0[(17792+col+1)*16-1-:16];
                next_layer_0[4479-:16] = layer_0[4479-:16] + layer_input[4479-:16]*kernel_0[(17856+col+1)*16-1-:16];
                next_layer_0[4495-:16] = layer_0[4495-:16] + layer_input[4495-:16]*kernel_0[(17920+col+1)*16-1-:16];
                next_layer_0[4511-:16] = layer_0[4511-:16] + layer_input[4511-:16]*kernel_0[(17984+col+1)*16-1-:16];
                next_layer_0[4527-:16] = layer_0[4527-:16] + layer_input[4527-:16]*kernel_0[(18048+col+1)*16-1-:16];
                next_layer_0[4543-:16] = layer_0[4543-:16] + layer_input[4543-:16]*kernel_0[(18112+col+1)*16-1-:16];
                next_layer_0[4559-:16] = layer_0[4559-:16] + layer_input[4559-:16]*kernel_0[(18176+col+1)*16-1-:16];
                next_layer_0[4575-:16] = layer_0[4575-:16] + layer_input[4575-:16]*kernel_0[(18240+col+1)*16-1-:16];
                next_layer_0[4591-:16] = layer_0[4591-:16] + layer_input[4591-:16]*kernel_0[(18304+col+1)*16-1-:16];
                next_layer_0[4607-:16] = layer_0[4607-:16] + layer_input[4607-:16]*kernel_0[(18368+col+1)*16-1-:16];
                next_layer_0[4623-:16] = layer_0[4623-:16] + layer_input[4623-:16]*kernel_0[(18432+col+1)*16-1-:16];
                next_layer_0[4639-:16] = layer_0[4639-:16] + layer_input[4639-:16]*kernel_0[(18496+col+1)*16-1-:16];
                next_layer_0[4655-:16] = layer_0[4655-:16] + layer_input[4655-:16]*kernel_0[(18560+col+1)*16-1-:16];
                next_layer_0[4671-:16] = layer_0[4671-:16] + layer_input[4671-:16]*kernel_0[(18624+col+1)*16-1-:16];
                next_layer_0[4687-:16] = layer_0[4687-:16] + layer_input[4687-:16]*kernel_0[(18688+col+1)*16-1-:16];
                next_layer_0[4703-:16] = layer_0[4703-:16] + layer_input[4703-:16]*kernel_0[(18752+col+1)*16-1-:16];
                next_layer_0[4719-:16] = layer_0[4719-:16] + layer_input[4719-:16]*kernel_0[(18816+col+1)*16-1-:16];
                next_layer_0[4735-:16] = layer_0[4735-:16] + layer_input[4735-:16]*kernel_0[(18880+col+1)*16-1-:16];
                next_layer_0[4751-:16] = layer_0[4751-:16] + layer_input[4751-:16]*kernel_0[(18944+col+1)*16-1-:16];
                next_layer_0[4767-:16] = layer_0[4767-:16] + layer_input[4767-:16]*kernel_0[(19008+col+1)*16-1-:16];
                next_layer_0[4783-:16] = layer_0[4783-:16] + layer_input[4783-:16]*kernel_0[(19072+col+1)*16-1-:16];
                next_layer_0[4799-:16] = layer_0[4799-:16] + layer_input[4799-:16]*kernel_0[(19136+col+1)*16-1-:16];
                next_layer_0[4815-:16] = layer_0[4815-:16] + layer_input[4815-:16]*kernel_0[(19200+col+1)*16-1-:16];
                next_layer_0[4831-:16] = layer_0[4831-:16] + layer_input[4831-:16]*kernel_0[(19264+col+1)*16-1-:16];
                next_layer_0[4847-:16] = layer_0[4847-:16] + layer_input[4847-:16]*kernel_0[(19328+col+1)*16-1-:16];
                next_layer_0[4863-:16] = layer_0[4863-:16] + layer_input[4863-:16]*kernel_0[(19392+col+1)*16-1-:16];
                next_layer_0[4879-:16] = layer_0[4879-:16] + layer_input[4879-:16]*kernel_0[(19456+col+1)*16-1-:16];
                next_layer_0[4895-:16] = layer_0[4895-:16] + layer_input[4895-:16]*kernel_0[(19520+col+1)*16-1-:16];
                next_layer_0[4911-:16] = layer_0[4911-:16] + layer_input[4911-:16]*kernel_0[(19584+col+1)*16-1-:16];
                next_layer_0[4927-:16] = layer_0[4927-:16] + layer_input[4927-:16]*kernel_0[(19648+col+1)*16-1-:16];
                next_layer_0[4943-:16] = layer_0[4943-:16] + layer_input[4943-:16]*kernel_0[(19712+col+1)*16-1-:16];
                next_layer_0[4959-:16] = layer_0[4959-:16] + layer_input[4959-:16]*kernel_0[(19776+col+1)*16-1-:16];
                next_layer_0[4975-:16] = layer_0[4975-:16] + layer_input[4975-:16]*kernel_0[(19840+col+1)*16-1-:16];
                next_layer_0[4991-:16] = layer_0[4991-:16] + layer_input[4991-:16]*kernel_0[(19904+col+1)*16-1-:16];
                next_layer_0[5007-:16] = layer_0[5007-:16] + layer_input[5007-:16]*kernel_0[(19968+col+1)*16-1-:16];
                next_layer_0[5023-:16] = layer_0[5023-:16] + layer_input[5023-:16]*kernel_0[(20032+col+1)*16-1-:16];
                next_layer_0[5039-:16] = layer_0[5039-:16] + layer_input[5039-:16]*kernel_0[(20096+col+1)*16-1-:16];
                next_layer_0[5055-:16] = layer_0[5055-:16] + layer_input[5055-:16]*kernel_0[(20160+col+1)*16-1-:16];
                next_layer_0[5071-:16] = layer_0[5071-:16] + layer_input[5071-:16]*kernel_0[(20224+col+1)*16-1-:16];
                next_layer_0[5087-:16] = layer_0[5087-:16] + layer_input[5087-:16]*kernel_0[(20288+col+1)*16-1-:16];
                next_layer_0[5103-:16] = layer_0[5103-:16] + layer_input[5103-:16]*kernel_0[(20352+col+1)*16-1-:16];
                next_layer_0[5119-:16] = layer_0[5119-:16] + layer_input[5119-:16]*kernel_0[(20416+col+1)*16-1-:16];
                next_layer_0[5135-:16] = layer_0[5135-:16] + layer_input[5135-:16]*kernel_0[(20480+col+1)*16-1-:16];
                next_layer_0[5151-:16] = layer_0[5151-:16] + layer_input[5151-:16]*kernel_0[(20544+col+1)*16-1-:16];
                next_layer_0[5167-:16] = layer_0[5167-:16] + layer_input[5167-:16]*kernel_0[(20608+col+1)*16-1-:16];
                next_layer_0[5183-:16] = layer_0[5183-:16] + layer_input[5183-:16]*kernel_0[(20672+col+1)*16-1-:16];
                next_layer_0[5199-:16] = layer_0[5199-:16] + layer_input[5199-:16]*kernel_0[(20736+col+1)*16-1-:16];
                next_layer_0[5215-:16] = layer_0[5215-:16] + layer_input[5215-:16]*kernel_0[(20800+col+1)*16-1-:16];
                next_layer_0[5231-:16] = layer_0[5231-:16] + layer_input[5231-:16]*kernel_0[(20864+col+1)*16-1-:16];
                next_layer_0[5247-:16] = layer_0[5247-:16] + layer_input[5247-:16]*kernel_0[(20928+col+1)*16-1-:16];
                next_layer_0[5263-:16] = layer_0[5263-:16] + layer_input[5263-:16]*kernel_0[(20992+col+1)*16-1-:16];
                next_layer_0[5279-:16] = layer_0[5279-:16] + layer_input[5279-:16]*kernel_0[(21056+col+1)*16-1-:16];
                next_layer_0[5295-:16] = layer_0[5295-:16] + layer_input[5295-:16]*kernel_0[(21120+col+1)*16-1-:16];
                next_layer_0[5311-:16] = layer_0[5311-:16] + layer_input[5311-:16]*kernel_0[(21184+col+1)*16-1-:16];
                next_layer_0[5327-:16] = layer_0[5327-:16] + layer_input[5327-:16]*kernel_0[(21248+col+1)*16-1-:16];
                next_layer_0[5343-:16] = layer_0[5343-:16] + layer_input[5343-:16]*kernel_0[(21312+col+1)*16-1-:16];
                next_layer_0[5359-:16] = layer_0[5359-:16] + layer_input[5359-:16]*kernel_0[(21376+col+1)*16-1-:16];
                next_layer_0[5375-:16] = layer_0[5375-:16] + layer_input[5375-:16]*kernel_0[(21440+col+1)*16-1-:16];
                next_layer_0[5391-:16] = layer_0[5391-:16] + layer_input[5391-:16]*kernel_0[(21504+col+1)*16-1-:16];
                next_layer_0[5407-:16] = layer_0[5407-:16] + layer_input[5407-:16]*kernel_0[(21568+col+1)*16-1-:16];
                next_layer_0[5423-:16] = layer_0[5423-:16] + layer_input[5423-:16]*kernel_0[(21632+col+1)*16-1-:16];
                next_layer_0[5439-:16] = layer_0[5439-:16] + layer_input[5439-:16]*kernel_0[(21696+col+1)*16-1-:16];
                next_layer_0[5455-:16] = layer_0[5455-:16] + layer_input[5455-:16]*kernel_0[(21760+col+1)*16-1-:16];
                next_layer_0[5471-:16] = layer_0[5471-:16] + layer_input[5471-:16]*kernel_0[(21824+col+1)*16-1-:16];
                next_layer_0[5487-:16] = layer_0[5487-:16] + layer_input[5487-:16]*kernel_0[(21888+col+1)*16-1-:16];
                next_layer_0[5503-:16] = layer_0[5503-:16] + layer_input[5503-:16]*kernel_0[(21952+col+1)*16-1-:16];
                next_layer_0[5519-:16] = layer_0[5519-:16] + layer_input[5519-:16]*kernel_0[(22016+col+1)*16-1-:16];
                next_layer_0[5535-:16] = layer_0[5535-:16] + layer_input[5535-:16]*kernel_0[(22080+col+1)*16-1-:16];
                next_layer_0[5551-:16] = layer_0[5551-:16] + layer_input[5551-:16]*kernel_0[(22144+col+1)*16-1-:16];
                next_layer_0[5567-:16] = layer_0[5567-:16] + layer_input[5567-:16]*kernel_0[(22208+col+1)*16-1-:16];
                next_layer_0[5583-:16] = layer_0[5583-:16] + layer_input[5583-:16]*kernel_0[(22272+col+1)*16-1-:16];
                next_layer_0[5599-:16] = layer_0[5599-:16] + layer_input[5599-:16]*kernel_0[(22336+col+1)*16-1-:16];
                next_layer_0[5615-:16] = layer_0[5615-:16] + layer_input[5615-:16]*kernel_0[(22400+col+1)*16-1-:16];
                next_layer_0[5631-:16] = layer_0[5631-:16] + layer_input[5631-:16]*kernel_0[(22464+col+1)*16-1-:16];
                next_layer_0[5647-:16] = layer_0[5647-:16] + layer_input[5647-:16]*kernel_0[(22528+col+1)*16-1-:16];
                next_layer_0[5663-:16] = layer_0[5663-:16] + layer_input[5663-:16]*kernel_0[(22592+col+1)*16-1-:16];
                next_layer_0[5679-:16] = layer_0[5679-:16] + layer_input[5679-:16]*kernel_0[(22656+col+1)*16-1-:16];
                next_layer_0[5695-:16] = layer_0[5695-:16] + layer_input[5695-:16]*kernel_0[(22720+col+1)*16-1-:16];
                next_layer_0[5711-:16] = layer_0[5711-:16] + layer_input[5711-:16]*kernel_0[(22784+col+1)*16-1-:16];
                next_layer_0[5727-:16] = layer_0[5727-:16] + layer_input[5727-:16]*kernel_0[(22848+col+1)*16-1-:16];
                next_layer_0[5743-:16] = layer_0[5743-:16] + layer_input[5743-:16]*kernel_0[(22912+col+1)*16-1-:16];
                next_layer_0[5759-:16] = layer_0[5759-:16] + layer_input[5759-:16]*kernel_0[(22976+col+1)*16-1-:16];
                next_layer_0[5775-:16] = layer_0[5775-:16] + layer_input[5775-:16]*kernel_0[(23040+col+1)*16-1-:16];
                next_layer_0[5791-:16] = layer_0[5791-:16] + layer_input[5791-:16]*kernel_0[(23104+col+1)*16-1-:16];
                next_layer_0[5807-:16] = layer_0[5807-:16] + layer_input[5807-:16]*kernel_0[(23168+col+1)*16-1-:16];
                next_layer_0[5823-:16] = layer_0[5823-:16] + layer_input[5823-:16]*kernel_0[(23232+col+1)*16-1-:16];
                next_layer_0[5839-:16] = layer_0[5839-:16] + layer_input[5839-:16]*kernel_0[(23296+col+1)*16-1-:16];
                next_layer_0[5855-:16] = layer_0[5855-:16] + layer_input[5855-:16]*kernel_0[(23360+col+1)*16-1-:16];
                next_layer_0[5871-:16] = layer_0[5871-:16] + layer_input[5871-:16]*kernel_0[(23424+col+1)*16-1-:16];
                next_layer_0[5887-:16] = layer_0[5887-:16] + layer_input[5887-:16]*kernel_0[(23488+col+1)*16-1-:16];
                next_layer_0[5903-:16] = layer_0[5903-:16] + layer_input[5903-:16]*kernel_0[(23552+col+1)*16-1-:16];
                next_layer_0[5919-:16] = layer_0[5919-:16] + layer_input[5919-:16]*kernel_0[(23616+col+1)*16-1-:16];
                next_layer_0[5935-:16] = layer_0[5935-:16] + layer_input[5935-:16]*kernel_0[(23680+col+1)*16-1-:16];
                next_layer_0[5951-:16] = layer_0[5951-:16] + layer_input[5951-:16]*kernel_0[(23744+col+1)*16-1-:16];
                next_layer_0[5967-:16] = layer_0[5967-:16] + layer_input[5967-:16]*kernel_0[(23808+col+1)*16-1-:16];
                next_layer_0[5983-:16] = layer_0[5983-:16] + layer_input[5983-:16]*kernel_0[(23872+col+1)*16-1-:16];
                next_layer_0[5999-:16] = layer_0[5999-:16] + layer_input[5999-:16]*kernel_0[(23936+col+1)*16-1-:16];
                next_layer_0[6015-:16] = layer_0[6015-:16] + layer_input[6015-:16]*kernel_0[(24000+col+1)*16-1-:16];
                next_layer_0[6031-:16] = layer_0[6031-:16] + layer_input[6031-:16]*kernel_0[(24064+col+1)*16-1-:16];
                next_layer_0[6047-:16] = layer_0[6047-:16] + layer_input[6047-:16]*kernel_0[(24128+col+1)*16-1-:16];
                next_layer_0[6063-:16] = layer_0[6063-:16] + layer_input[6063-:16]*kernel_0[(24192+col+1)*16-1-:16];
                next_layer_0[6079-:16] = layer_0[6079-:16] + layer_input[6079-:16]*kernel_0[(24256+col+1)*16-1-:16];
                next_layer_0[6095-:16] = layer_0[6095-:16] + layer_input[6095-:16]*kernel_0[(24320+col+1)*16-1-:16];
                next_layer_0[6111-:16] = layer_0[6111-:16] + layer_input[6111-:16]*kernel_0[(24384+col+1)*16-1-:16];
                next_layer_0[6127-:16] = layer_0[6127-:16] + layer_input[6127-:16]*kernel_0[(24448+col+1)*16-1-:16];
                next_layer_0[6143-:16] = layer_0[6143-:16] + layer_input[6143-:16]*kernel_0[(24512+col+1)*16-1-:16];
                next_layer_0[6159-:16] = layer_0[6159-:16] + layer_input[6159-:16]*kernel_0[(24576+col+1)*16-1-:16];
                next_layer_0[6175-:16] = layer_0[6175-:16] + layer_input[6175-:16]*kernel_0[(24640+col+1)*16-1-:16];
                next_layer_0[6191-:16] = layer_0[6191-:16] + layer_input[6191-:16]*kernel_0[(24704+col+1)*16-1-:16];
                next_layer_0[6207-:16] = layer_0[6207-:16] + layer_input[6207-:16]*kernel_0[(24768+col+1)*16-1-:16];
                next_layer_0[6223-:16] = layer_0[6223-:16] + layer_input[6223-:16]*kernel_0[(24832+col+1)*16-1-:16];
                next_layer_0[6239-:16] = layer_0[6239-:16] + layer_input[6239-:16]*kernel_0[(24896+col+1)*16-1-:16];
                next_layer_0[6255-:16] = layer_0[6255-:16] + layer_input[6255-:16]*kernel_0[(24960+col+1)*16-1-:16];
                next_layer_0[6271-:16] = layer_0[6271-:16] + layer_input[6271-:16]*kernel_0[(25024+col+1)*16-1-:16];
                next_layer_0[6287-:16] = layer_0[6287-:16] + layer_input[6287-:16]*kernel_0[(25088+col+1)*16-1-:16];
                next_layer_0[6303-:16] = layer_0[6303-:16] + layer_input[6303-:16]*kernel_0[(25152+col+1)*16-1-:16];
                next_layer_0[6319-:16] = layer_0[6319-:16] + layer_input[6319-:16]*kernel_0[(25216+col+1)*16-1-:16];
                next_layer_0[6335-:16] = layer_0[6335-:16] + layer_input[6335-:16]*kernel_0[(25280+col+1)*16-1-:16];
                next_layer_0[6351-:16] = layer_0[6351-:16] + layer_input[6351-:16]*kernel_0[(25344+col+1)*16-1-:16];
                next_layer_0[6367-:16] = layer_0[6367-:16] + layer_input[6367-:16]*kernel_0[(25408+col+1)*16-1-:16];
                next_layer_0[6383-:16] = layer_0[6383-:16] + layer_input[6383-:16]*kernel_0[(25472+col+1)*16-1-:16];
                next_layer_0[6399-:16] = layer_0[6399-:16] + layer_input[6399-:16]*kernel_0[(25536+col+1)*16-1-:16];
                next_layer_0[6415-:16] = layer_0[6415-:16] + layer_input[6415-:16]*kernel_0[(25600+col+1)*16-1-:16];
                next_layer_0[6431-:16] = layer_0[6431-:16] + layer_input[6431-:16]*kernel_0[(25664+col+1)*16-1-:16];
                next_layer_0[6447-:16] = layer_0[6447-:16] + layer_input[6447-:16]*kernel_0[(25728+col+1)*16-1-:16];
                next_layer_0[6463-:16] = layer_0[6463-:16] + layer_input[6463-:16]*kernel_0[(25792+col+1)*16-1-:16];
                next_layer_0[6479-:16] = layer_0[6479-:16] + layer_input[6479-:16]*kernel_0[(25856+col+1)*16-1-:16];
                next_layer_0[6495-:16] = layer_0[6495-:16] + layer_input[6495-:16]*kernel_0[(25920+col+1)*16-1-:16];
                next_layer_0[6511-:16] = layer_0[6511-:16] + layer_input[6511-:16]*kernel_0[(25984+col+1)*16-1-:16];
                next_layer_0[6527-:16] = layer_0[6527-:16] + layer_input[6527-:16]*kernel_0[(26048+col+1)*16-1-:16];
                next_layer_0[6543-:16] = layer_0[6543-:16] + layer_input[6543-:16]*kernel_0[(26112+col+1)*16-1-:16];
                next_layer_0[6559-:16] = layer_0[6559-:16] + layer_input[6559-:16]*kernel_0[(26176+col+1)*16-1-:16];
                next_layer_0[6575-:16] = layer_0[6575-:16] + layer_input[6575-:16]*kernel_0[(26240+col+1)*16-1-:16];
                next_layer_0[6591-:16] = layer_0[6591-:16] + layer_input[6591-:16]*kernel_0[(26304+col+1)*16-1-:16];
                next_layer_0[6607-:16] = layer_0[6607-:16] + layer_input[6607-:16]*kernel_0[(26368+col+1)*16-1-:16];
                next_layer_0[6623-:16] = layer_0[6623-:16] + layer_input[6623-:16]*kernel_0[(26432+col+1)*16-1-:16];
                next_layer_0[6639-:16] = layer_0[6639-:16] + layer_input[6639-:16]*kernel_0[(26496+col+1)*16-1-:16];
                next_layer_0[6655-:16] = layer_0[6655-:16] + layer_input[6655-:16]*kernel_0[(26560+col+1)*16-1-:16];
                next_layer_0[6671-:16] = layer_0[6671-:16] + layer_input[6671-:16]*kernel_0[(26624+col+1)*16-1-:16];
                next_layer_0[6687-:16] = layer_0[6687-:16] + layer_input[6687-:16]*kernel_0[(26688+col+1)*16-1-:16];
                next_layer_0[6703-:16] = layer_0[6703-:16] + layer_input[6703-:16]*kernel_0[(26752+col+1)*16-1-:16];
                next_layer_0[6719-:16] = layer_0[6719-:16] + layer_input[6719-:16]*kernel_0[(26816+col+1)*16-1-:16];
                next_layer_0[6735-:16] = layer_0[6735-:16] + layer_input[6735-:16]*kernel_0[(26880+col+1)*16-1-:16];
                next_layer_0[6751-:16] = layer_0[6751-:16] + layer_input[6751-:16]*kernel_0[(26944+col+1)*16-1-:16];
                next_layer_0[6767-:16] = layer_0[6767-:16] + layer_input[6767-:16]*kernel_0[(27008+col+1)*16-1-:16];
                next_layer_0[6783-:16] = layer_0[6783-:16] + layer_input[6783-:16]*kernel_0[(27072+col+1)*16-1-:16];
                next_layer_0[6799-:16] = layer_0[6799-:16] + layer_input[6799-:16]*kernel_0[(27136+col+1)*16-1-:16];
                next_layer_0[6815-:16] = layer_0[6815-:16] + layer_input[6815-:16]*kernel_0[(27200+col+1)*16-1-:16];
                next_layer_0[6831-:16] = layer_0[6831-:16] + layer_input[6831-:16]*kernel_0[(27264+col+1)*16-1-:16];
                next_layer_0[6847-:16] = layer_0[6847-:16] + layer_input[6847-:16]*kernel_0[(27328+col+1)*16-1-:16];
                next_layer_0[6863-:16] = layer_0[6863-:16] + layer_input[6863-:16]*kernel_0[(27392+col+1)*16-1-:16];
                next_layer_0[6879-:16] = layer_0[6879-:16] + layer_input[6879-:16]*kernel_0[(27456+col+1)*16-1-:16];
                next_layer_0[6895-:16] = layer_0[6895-:16] + layer_input[6895-:16]*kernel_0[(27520+col+1)*16-1-:16];
                next_layer_0[6911-:16] = layer_0[6911-:16] + layer_input[6911-:16]*kernel_0[(27584+col+1)*16-1-:16];
                next_layer_0[6927-:16] = layer_0[6927-:16] + layer_input[6927-:16]*kernel_0[(27648+col+1)*16-1-:16];
                next_layer_0[6943-:16] = layer_0[6943-:16] + layer_input[6943-:16]*kernel_0[(27712+col+1)*16-1-:16];
                next_layer_0[6959-:16] = layer_0[6959-:16] + layer_input[6959-:16]*kernel_0[(27776+col+1)*16-1-:16];
                next_layer_0[6975-:16] = layer_0[6975-:16] + layer_input[6975-:16]*kernel_0[(27840+col+1)*16-1-:16];
                next_layer_0[6991-:16] = layer_0[6991-:16] + layer_input[6991-:16]*kernel_0[(27904+col+1)*16-1-:16];
                next_layer_0[7007-:16] = layer_0[7007-:16] + layer_input[7007-:16]*kernel_0[(27968+col+1)*16-1-:16];
                next_layer_0[7023-:16] = layer_0[7023-:16] + layer_input[7023-:16]*kernel_0[(28032+col+1)*16-1-:16];
                next_layer_0[7039-:16] = layer_0[7039-:16] + layer_input[7039-:16]*kernel_0[(28096+col+1)*16-1-:16];
                next_layer_0[7055-:16] = layer_0[7055-:16] + layer_input[7055-:16]*kernel_0[(28160+col+1)*16-1-:16];
                next_layer_0[7071-:16] = layer_0[7071-:16] + layer_input[7071-:16]*kernel_0[(28224+col+1)*16-1-:16];
                next_layer_0[7087-:16] = layer_0[7087-:16] + layer_input[7087-:16]*kernel_0[(28288+col+1)*16-1-:16];
                next_layer_0[7103-:16] = layer_0[7103-:16] + layer_input[7103-:16]*kernel_0[(28352+col+1)*16-1-:16];
                next_layer_0[7119-:16] = layer_0[7119-:16] + layer_input[7119-:16]*kernel_0[(28416+col+1)*16-1-:16];
                next_layer_0[7135-:16] = layer_0[7135-:16] + layer_input[7135-:16]*kernel_0[(28480+col+1)*16-1-:16];
                next_layer_0[7151-:16] = layer_0[7151-:16] + layer_input[7151-:16]*kernel_0[(28544+col+1)*16-1-:16];
                next_layer_0[7167-:16] = layer_0[7167-:16] + layer_input[7167-:16]*kernel_0[(28608+col+1)*16-1-:16];
                next_layer_0[7183-:16] = layer_0[7183-:16] + layer_input[7183-:16]*kernel_0[(28672+col+1)*16-1-:16];
                next_layer_0[7199-:16] = layer_0[7199-:16] + layer_input[7199-:16]*kernel_0[(28736+col+1)*16-1-:16];
                next_layer_0[7215-:16] = layer_0[7215-:16] + layer_input[7215-:16]*kernel_0[(28800+col+1)*16-1-:16];
                next_layer_0[7231-:16] = layer_0[7231-:16] + layer_input[7231-:16]*kernel_0[(28864+col+1)*16-1-:16];
                next_layer_0[7247-:16] = layer_0[7247-:16] + layer_input[7247-:16]*kernel_0[(28928+col+1)*16-1-:16];
                next_layer_0[7263-:16] = layer_0[7263-:16] + layer_input[7263-:16]*kernel_0[(28992+col+1)*16-1-:16];
                next_layer_0[7279-:16] = layer_0[7279-:16] + layer_input[7279-:16]*kernel_0[(29056+col+1)*16-1-:16];
                next_layer_0[7295-:16] = layer_0[7295-:16] + layer_input[7295-:16]*kernel_0[(29120+col+1)*16-1-:16];
                next_layer_0[7311-:16] = layer_0[7311-:16] + layer_input[7311-:16]*kernel_0[(29184+col+1)*16-1-:16];
                next_layer_0[7327-:16] = layer_0[7327-:16] + layer_input[7327-:16]*kernel_0[(29248+col+1)*16-1-:16];
                next_layer_0[7343-:16] = layer_0[7343-:16] + layer_input[7343-:16]*kernel_0[(29312+col+1)*16-1-:16];
                next_layer_0[7359-:16] = layer_0[7359-:16] + layer_input[7359-:16]*kernel_0[(29376+col+1)*16-1-:16];
                next_layer_0[7375-:16] = layer_0[7375-:16] + layer_input[7375-:16]*kernel_0[(29440+col+1)*16-1-:16];
                next_layer_0[7391-:16] = layer_0[7391-:16] + layer_input[7391-:16]*kernel_0[(29504+col+1)*16-1-:16];
                next_layer_0[7407-:16] = layer_0[7407-:16] + layer_input[7407-:16]*kernel_0[(29568+col+1)*16-1-:16];
                next_layer_0[7423-:16] = layer_0[7423-:16] + layer_input[7423-:16]*kernel_0[(29632+col+1)*16-1-:16];
                next_layer_0[7439-:16] = layer_0[7439-:16] + layer_input[7439-:16]*kernel_0[(29696+col+1)*16-1-:16];
                next_layer_0[7455-:16] = layer_0[7455-:16] + layer_input[7455-:16]*kernel_0[(29760+col+1)*16-1-:16];
                next_layer_0[7471-:16] = layer_0[7471-:16] + layer_input[7471-:16]*kernel_0[(29824+col+1)*16-1-:16];
                next_layer_0[7487-:16] = layer_0[7487-:16] + layer_input[7487-:16]*kernel_0[(29888+col+1)*16-1-:16];
                next_layer_0[7503-:16] = layer_0[7503-:16] + layer_input[7503-:16]*kernel_0[(29952+col+1)*16-1-:16];
                next_layer_0[7519-:16] = layer_0[7519-:16] + layer_input[7519-:16]*kernel_0[(30016+col+1)*16-1-:16];
                next_layer_0[7535-:16] = layer_0[7535-:16] + layer_input[7535-:16]*kernel_0[(30080+col+1)*16-1-:16];
                next_layer_0[7551-:16] = layer_0[7551-:16] + layer_input[7551-:16]*kernel_0[(30144+col+1)*16-1-:16];
                next_layer_0[7567-:16] = layer_0[7567-:16] + layer_input[7567-:16]*kernel_0[(30208+col+1)*16-1-:16];
                next_layer_0[7583-:16] = layer_0[7583-:16] + layer_input[7583-:16]*kernel_0[(30272+col+1)*16-1-:16];
                next_layer_0[7599-:16] = layer_0[7599-:16] + layer_input[7599-:16]*kernel_0[(30336+col+1)*16-1-:16];
                next_layer_0[7615-:16] = layer_0[7615-:16] + layer_input[7615-:16]*kernel_0[(30400+col+1)*16-1-:16];
                next_layer_0[7631-:16] = layer_0[7631-:16] + layer_input[7631-:16]*kernel_0[(30464+col+1)*16-1-:16];
                next_layer_0[7647-:16] = layer_0[7647-:16] + layer_input[7647-:16]*kernel_0[(30528+col+1)*16-1-:16];
                next_layer_0[7663-:16] = layer_0[7663-:16] + layer_input[7663-:16]*kernel_0[(30592+col+1)*16-1-:16];
                next_layer_0[7679-:16] = layer_0[7679-:16] + layer_input[7679-:16]*kernel_0[(30656+col+1)*16-1-:16];
                next_layer_0[7695-:16] = layer_0[7695-:16] + layer_input[7695-:16]*kernel_0[(30720+col+1)*16-1-:16];
                next_layer_0[7711-:16] = layer_0[7711-:16] + layer_input[7711-:16]*kernel_0[(30784+col+1)*16-1-:16];
                next_layer_0[7727-:16] = layer_0[7727-:16] + layer_input[7727-:16]*kernel_0[(30848+col+1)*16-1-:16];
                next_layer_0[7743-:16] = layer_0[7743-:16] + layer_input[7743-:16]*kernel_0[(30912+col+1)*16-1-:16];
                next_layer_0[7759-:16] = layer_0[7759-:16] + layer_input[7759-:16]*kernel_0[(30976+col+1)*16-1-:16];
                next_layer_0[7775-:16] = layer_0[7775-:16] + layer_input[7775-:16]*kernel_0[(31040+col+1)*16-1-:16];
                next_layer_0[7791-:16] = layer_0[7791-:16] + layer_input[7791-:16]*kernel_0[(31104+col+1)*16-1-:16];
                next_layer_0[7807-:16] = layer_0[7807-:16] + layer_input[7807-:16]*kernel_0[(31168+col+1)*16-1-:16];
                next_layer_0[7823-:16] = layer_0[7823-:16] + layer_input[7823-:16]*kernel_0[(31232+col+1)*16-1-:16];
                next_layer_0[7839-:16] = layer_0[7839-:16] + layer_input[7839-:16]*kernel_0[(31296+col+1)*16-1-:16];
                next_layer_0[7855-:16] = layer_0[7855-:16] + layer_input[7855-:16]*kernel_0[(31360+col+1)*16-1-:16];
                next_layer_0[7871-:16] = layer_0[7871-:16] + layer_input[7871-:16]*kernel_0[(31424+col+1)*16-1-:16];
                next_layer_0[7887-:16] = layer_0[7887-:16] + layer_input[7887-:16]*kernel_0[(31488+col+1)*16-1-:16];
                next_layer_0[7903-:16] = layer_0[7903-:16] + layer_input[7903-:16]*kernel_0[(31552+col+1)*16-1-:16];
                next_layer_0[7919-:16] = layer_0[7919-:16] + layer_input[7919-:16]*kernel_0[(31616+col+1)*16-1-:16];
                next_layer_0[7935-:16] = layer_0[7935-:16] + layer_input[7935-:16]*kernel_0[(31680+col+1)*16-1-:16];
                next_layer_0[7951-:16] = layer_0[7951-:16] + layer_input[7951-:16]*kernel_0[(31744+col+1)*16-1-:16];
                next_layer_0[7967-:16] = layer_0[7967-:16] + layer_input[7967-:16]*kernel_0[(31808+col+1)*16-1-:16];
                next_layer_0[7983-:16] = layer_0[7983-:16] + layer_input[7983-:16]*kernel_0[(31872+col+1)*16-1-:16];
                next_layer_0[7999-:16] = layer_0[7999-:16] + layer_input[7999-:16]*kernel_0[(31936+col+1)*16-1-:16];
                next_layer_0[8015-:16] = layer_0[8015-:16] + layer_input[8015-:16]*kernel_0[(32000+col+1)*16-1-:16];
                next_layer_0[8031-:16] = layer_0[8031-:16] + layer_input[8031-:16]*kernel_0[(32064+col+1)*16-1-:16];
                next_layer_0[8047-:16] = layer_0[8047-:16] + layer_input[8047-:16]*kernel_0[(32128+col+1)*16-1-:16];
                next_layer_0[8063-:16] = layer_0[8063-:16] + layer_input[8063-:16]*kernel_0[(32192+col+1)*16-1-:16];
                next_layer_0[8079-:16] = layer_0[8079-:16] + layer_input[8079-:16]*kernel_0[(32256+col+1)*16-1-:16];
                next_layer_0[8095-:16] = layer_0[8095-:16] + layer_input[8095-:16]*kernel_0[(32320+col+1)*16-1-:16];
                next_layer_0[8111-:16] = layer_0[8111-:16] + layer_input[8111-:16]*kernel_0[(32384+col+1)*16-1-:16];
                next_layer_0[8127-:16] = layer_0[8127-:16] + layer_input[8127-:16]*kernel_0[(32448+col+1)*16-1-:16];
                next_layer_0[8143-:16] = layer_0[8143-:16] + layer_input[8143-:16]*kernel_0[(32512+col+1)*16-1-:16];
                next_layer_0[8159-:16] = layer_0[8159-:16] + layer_input[8159-:16]*kernel_0[(32576+col+1)*16-1-:16];
                next_layer_0[8175-:16] = layer_0[8175-:16] + layer_input[8175-:16]*kernel_0[(32640+col+1)*16-1-:16];
                next_layer_0[8191-:16] = layer_0[8191-:16] + layer_input[8191-:16]*kernel_0[(32704+col+1)*16-1-:16];
                next_layer_0[8207-:16] = layer_0[8207-:16] + layer_input[8207-:16]*kernel_0[(32768+col+1)*16-1-:16];
                next_layer_0[8223-:16] = layer_0[8223-:16] + layer_input[8223-:16]*kernel_0[(32832+col+1)*16-1-:16];
                next_layer_0[8239-:16] = layer_0[8239-:16] + layer_input[8239-:16]*kernel_0[(32896+col+1)*16-1-:16];
                next_layer_0[8255-:16] = layer_0[8255-:16] + layer_input[8255-:16]*kernel_0[(32960+col+1)*16-1-:16];
                next_layer_0[8271-:16] = layer_0[8271-:16] + layer_input[8271-:16]*kernel_0[(33024+col+1)*16-1-:16];
                next_layer_0[8287-:16] = layer_0[8287-:16] + layer_input[8287-:16]*kernel_0[(33088+col+1)*16-1-:16];
                next_layer_0[8303-:16] = layer_0[8303-:16] + layer_input[8303-:16]*kernel_0[(33152+col+1)*16-1-:16];
                next_layer_0[8319-:16] = layer_0[8319-:16] + layer_input[8319-:16]*kernel_0[(33216+col+1)*16-1-:16];
                next_layer_0[8335-:16] = layer_0[8335-:16] + layer_input[8335-:16]*kernel_0[(33280+col+1)*16-1-:16];
                next_layer_0[8351-:16] = layer_0[8351-:16] + layer_input[8351-:16]*kernel_0[(33344+col+1)*16-1-:16];
                next_layer_0[8367-:16] = layer_0[8367-:16] + layer_input[8367-:16]*kernel_0[(33408+col+1)*16-1-:16];
                next_layer_0[8383-:16] = layer_0[8383-:16] + layer_input[8383-:16]*kernel_0[(33472+col+1)*16-1-:16];
                next_layer_0[8399-:16] = layer_0[8399-:16] + layer_input[8399-:16]*kernel_0[(33536+col+1)*16-1-:16];
                next_layer_0[8415-:16] = layer_0[8415-:16] + layer_input[8415-:16]*kernel_0[(33600+col+1)*16-1-:16];
                next_layer_0[8431-:16] = layer_0[8431-:16] + layer_input[8431-:16]*kernel_0[(33664+col+1)*16-1-:16];
                next_layer_0[8447-:16] = layer_0[8447-:16] + layer_input[8447-:16]*kernel_0[(33728+col+1)*16-1-:16];
                next_layer_0[8463-:16] = layer_0[8463-:16] + layer_input[8463-:16]*kernel_0[(33792+col+1)*16-1-:16];
                next_layer_0[8479-:16] = layer_0[8479-:16] + layer_input[8479-:16]*kernel_0[(33856+col+1)*16-1-:16];
                next_layer_0[8495-:16] = layer_0[8495-:16] + layer_input[8495-:16]*kernel_0[(33920+col+1)*16-1-:16];
                next_layer_0[8511-:16] = layer_0[8511-:16] + layer_input[8511-:16]*kernel_0[(33984+col+1)*16-1-:16];
                next_layer_0[8527-:16] = layer_0[8527-:16] + layer_input[8527-:16]*kernel_0[(34048+col+1)*16-1-:16];
                next_layer_0[8543-:16] = layer_0[8543-:16] + layer_input[8543-:16]*kernel_0[(34112+col+1)*16-1-:16];
                next_layer_0[8559-:16] = layer_0[8559-:16] + layer_input[8559-:16]*kernel_0[(34176+col+1)*16-1-:16];
                next_layer_0[8575-:16] = layer_0[8575-:16] + layer_input[8575-:16]*kernel_0[(34240+col+1)*16-1-:16];
                next_layer_0[8591-:16] = layer_0[8591-:16] + layer_input[8591-:16]*kernel_0[(34304+col+1)*16-1-:16];
                next_layer_0[8607-:16] = layer_0[8607-:16] + layer_input[8607-:16]*kernel_0[(34368+col+1)*16-1-:16];
                next_layer_0[8623-:16] = layer_0[8623-:16] + layer_input[8623-:16]*kernel_0[(34432+col+1)*16-1-:16];
                next_layer_0[8639-:16] = layer_0[8639-:16] + layer_input[8639-:16]*kernel_0[(34496+col+1)*16-1-:16];
                next_layer_0[8655-:16] = layer_0[8655-:16] + layer_input[8655-:16]*kernel_0[(34560+col+1)*16-1-:16];
                next_layer_0[8671-:16] = layer_0[8671-:16] + layer_input[8671-:16]*kernel_0[(34624+col+1)*16-1-:16];
                next_layer_0[8687-:16] = layer_0[8687-:16] + layer_input[8687-:16]*kernel_0[(34688+col+1)*16-1-:16];
                next_layer_0[8703-:16] = layer_0[8703-:16] + layer_input[8703-:16]*kernel_0[(34752+col+1)*16-1-:16];
                next_layer_0[8719-:16] = layer_0[8719-:16] + layer_input[8719-:16]*kernel_0[(34816+col+1)*16-1-:16];
                next_layer_0[8735-:16] = layer_0[8735-:16] + layer_input[8735-:16]*kernel_0[(34880+col+1)*16-1-:16];
                next_layer_0[8751-:16] = layer_0[8751-:16] + layer_input[8751-:16]*kernel_0[(34944+col+1)*16-1-:16];
                next_layer_0[8767-:16] = layer_0[8767-:16] + layer_input[8767-:16]*kernel_0[(35008+col+1)*16-1-:16];
                next_layer_0[8783-:16] = layer_0[8783-:16] + layer_input[8783-:16]*kernel_0[(35072+col+1)*16-1-:16];
                next_layer_0[8799-:16] = layer_0[8799-:16] + layer_input[8799-:16]*kernel_0[(35136+col+1)*16-1-:16];
                next_layer_0[8815-:16] = layer_0[8815-:16] + layer_input[8815-:16]*kernel_0[(35200+col+1)*16-1-:16];
                next_layer_0[8831-:16] = layer_0[8831-:16] + layer_input[8831-:16]*kernel_0[(35264+col+1)*16-1-:16];
                next_layer_0[8847-:16] = layer_0[8847-:16] + layer_input[8847-:16]*kernel_0[(35328+col+1)*16-1-:16];
                next_layer_0[8863-:16] = layer_0[8863-:16] + layer_input[8863-:16]*kernel_0[(35392+col+1)*16-1-:16];
                next_layer_0[8879-:16] = layer_0[8879-:16] + layer_input[8879-:16]*kernel_0[(35456+col+1)*16-1-:16];
                next_layer_0[8895-:16] = layer_0[8895-:16] + layer_input[8895-:16]*kernel_0[(35520+col+1)*16-1-:16];
                next_layer_0[8911-:16] = layer_0[8911-:16] + layer_input[8911-:16]*kernel_0[(35584+col+1)*16-1-:16];
                next_layer_0[8927-:16] = layer_0[8927-:16] + layer_input[8927-:16]*kernel_0[(35648+col+1)*16-1-:16];
                next_layer_0[8943-:16] = layer_0[8943-:16] + layer_input[8943-:16]*kernel_0[(35712+col+1)*16-1-:16];
                next_layer_0[8959-:16] = layer_0[8959-:16] + layer_input[8959-:16]*kernel_0[(35776+col+1)*16-1-:16];
                next_layer_0[8975-:16] = layer_0[8975-:16] + layer_input[8975-:16]*kernel_0[(35840+col+1)*16-1-:16];
                next_layer_0[8991-:16] = layer_0[8991-:16] + layer_input[8991-:16]*kernel_0[(35904+col+1)*16-1-:16];
                next_layer_0[9007-:16] = layer_0[9007-:16] + layer_input[9007-:16]*kernel_0[(35968+col+1)*16-1-:16];
                next_layer_0[9023-:16] = layer_0[9023-:16] + layer_input[9023-:16]*kernel_0[(36032+col+1)*16-1-:16];
                next_layer_0[9039-:16] = layer_0[9039-:16] + layer_input[9039-:16]*kernel_0[(36096+col+1)*16-1-:16];
                next_layer_0[9055-:16] = layer_0[9055-:16] + layer_input[9055-:16]*kernel_0[(36160+col+1)*16-1-:16];
                next_layer_0[9071-:16] = layer_0[9071-:16] + layer_input[9071-:16]*kernel_0[(36224+col+1)*16-1-:16];
                next_layer_0[9087-:16] = layer_0[9087-:16] + layer_input[9087-:16]*kernel_0[(36288+col+1)*16-1-:16];
                next_layer_0[9103-:16] = layer_0[9103-:16] + layer_input[9103-:16]*kernel_0[(36352+col+1)*16-1-:16];
                next_layer_0[9119-:16] = layer_0[9119-:16] + layer_input[9119-:16]*kernel_0[(36416+col+1)*16-1-:16];
                next_layer_0[9135-:16] = layer_0[9135-:16] + layer_input[9135-:16]*kernel_0[(36480+col+1)*16-1-:16];
                next_layer_0[9151-:16] = layer_0[9151-:16] + layer_input[9151-:16]*kernel_0[(36544+col+1)*16-1-:16];
                next_layer_0[9167-:16] = layer_0[9167-:16] + layer_input[9167-:16]*kernel_0[(36608+col+1)*16-1-:16];
                next_layer_0[9183-:16] = layer_0[9183-:16] + layer_input[9183-:16]*kernel_0[(36672+col+1)*16-1-:16];
                next_layer_0[9199-:16] = layer_0[9199-:16] + layer_input[9199-:16]*kernel_0[(36736+col+1)*16-1-:16];
                next_layer_0[9215-:16] = layer_0[9215-:16] + layer_input[9215-:16]*kernel_0[(36800+col+1)*16-1-:16];
                next_layer_0[9231-:16] = layer_0[9231-:16] + layer_input[9231-:16]*kernel_0[(36864+col+1)*16-1-:16];
                next_layer_0[9247-:16] = layer_0[9247-:16] + layer_input[9247-:16]*kernel_0[(36928+col+1)*16-1-:16];
                next_layer_0[9263-:16] = layer_0[9263-:16] + layer_input[9263-:16]*kernel_0[(36992+col+1)*16-1-:16];
                next_layer_0[9279-:16] = layer_0[9279-:16] + layer_input[9279-:16]*kernel_0[(37056+col+1)*16-1-:16];
                next_layer_0[9295-:16] = layer_0[9295-:16] + layer_input[9295-:16]*kernel_0[(37120+col+1)*16-1-:16];
                next_layer_0[9311-:16] = layer_0[9311-:16] + layer_input[9311-:16]*kernel_0[(37184+col+1)*16-1-:16];
                next_layer_0[9327-:16] = layer_0[9327-:16] + layer_input[9327-:16]*kernel_0[(37248+col+1)*16-1-:16];
                next_layer_0[9343-:16] = layer_0[9343-:16] + layer_input[9343-:16]*kernel_0[(37312+col+1)*16-1-:16];
                next_layer_0[9359-:16] = layer_0[9359-:16] + layer_input[9359-:16]*kernel_0[(37376+col+1)*16-1-:16];
                next_layer_0[9375-:16] = layer_0[9375-:16] + layer_input[9375-:16]*kernel_0[(37440+col+1)*16-1-:16];
                next_layer_0[9391-:16] = layer_0[9391-:16] + layer_input[9391-:16]*kernel_0[(37504+col+1)*16-1-:16];
                next_layer_0[9407-:16] = layer_0[9407-:16] + layer_input[9407-:16]*kernel_0[(37568+col+1)*16-1-:16];
                next_layer_0[9423-:16] = layer_0[9423-:16] + layer_input[9423-:16]*kernel_0[(37632+col+1)*16-1-:16];
                next_layer_0[9439-:16] = layer_0[9439-:16] + layer_input[9439-:16]*kernel_0[(37696+col+1)*16-1-:16];
                next_layer_0[9455-:16] = layer_0[9455-:16] + layer_input[9455-:16]*kernel_0[(37760+col+1)*16-1-:16];
                next_layer_0[9471-:16] = layer_0[9471-:16] + layer_input[9471-:16]*kernel_0[(37824+col+1)*16-1-:16];
                next_layer_0[9487-:16] = layer_0[9487-:16] + layer_input[9487-:16]*kernel_0[(37888+col+1)*16-1-:16];
                next_layer_0[9503-:16] = layer_0[9503-:16] + layer_input[9503-:16]*kernel_0[(37952+col+1)*16-1-:16];
                next_layer_0[9519-:16] = layer_0[9519-:16] + layer_input[9519-:16]*kernel_0[(38016+col+1)*16-1-:16];
                next_layer_0[9535-:16] = layer_0[9535-:16] + layer_input[9535-:16]*kernel_0[(38080+col+1)*16-1-:16];
                next_layer_0[9551-:16] = layer_0[9551-:16] + layer_input[9551-:16]*kernel_0[(38144+col+1)*16-1-:16];
                next_layer_0[9567-:16] = layer_0[9567-:16] + layer_input[9567-:16]*kernel_0[(38208+col+1)*16-1-:16];
                next_layer_0[9583-:16] = layer_0[9583-:16] + layer_input[9583-:16]*kernel_0[(38272+col+1)*16-1-:16];
                next_layer_0[9599-:16] = layer_0[9599-:16] + layer_input[9599-:16]*kernel_0[(38336+col+1)*16-1-:16];
                next_layer_0[9615-:16] = layer_0[9615-:16] + layer_input[9615-:16]*kernel_0[(38400+col+1)*16-1-:16];
                next_layer_0[9631-:16] = layer_0[9631-:16] + layer_input[9631-:16]*kernel_0[(38464+col+1)*16-1-:16];
                next_layer_0[9647-:16] = layer_0[9647-:16] + layer_input[9647-:16]*kernel_0[(38528+col+1)*16-1-:16];
                next_layer_0[9663-:16] = layer_0[9663-:16] + layer_input[9663-:16]*kernel_0[(38592+col+1)*16-1-:16];
                next_layer_0[9679-:16] = layer_0[9679-:16] + layer_input[9679-:16]*kernel_0[(38656+col+1)*16-1-:16];
                next_layer_0[9695-:16] = layer_0[9695-:16] + layer_input[9695-:16]*kernel_0[(38720+col+1)*16-1-:16];
                next_layer_0[9711-:16] = layer_0[9711-:16] + layer_input[9711-:16]*kernel_0[(38784+col+1)*16-1-:16];
                next_layer_0[9727-:16] = layer_0[9727-:16] + layer_input[9727-:16]*kernel_0[(38848+col+1)*16-1-:16];
                next_layer_0[9743-:16] = layer_0[9743-:16] + layer_input[9743-:16]*kernel_0[(38912+col+1)*16-1-:16];
                next_layer_0[9759-:16] = layer_0[9759-:16] + layer_input[9759-:16]*kernel_0[(38976+col+1)*16-1-:16];
                next_layer_0[9775-:16] = layer_0[9775-:16] + layer_input[9775-:16]*kernel_0[(39040+col+1)*16-1-:16];
                next_layer_0[9791-:16] = layer_0[9791-:16] + layer_input[9791-:16]*kernel_0[(39104+col+1)*16-1-:16];
                next_layer_0[9807-:16] = layer_0[9807-:16] + layer_input[9807-:16]*kernel_0[(39168+col+1)*16-1-:16];
                next_layer_0[9823-:16] = layer_0[9823-:16] + layer_input[9823-:16]*kernel_0[(39232+col+1)*16-1-:16];
                next_layer_0[9839-:16] = layer_0[9839-:16] + layer_input[9839-:16]*kernel_0[(39296+col+1)*16-1-:16];
                next_layer_0[9855-:16] = layer_0[9855-:16] + layer_input[9855-:16]*kernel_0[(39360+col+1)*16-1-:16];
                next_layer_0[9871-:16] = layer_0[9871-:16] + layer_input[9871-:16]*kernel_0[(39424+col+1)*16-1-:16];
                next_layer_0[9887-:16] = layer_0[9887-:16] + layer_input[9887-:16]*kernel_0[(39488+col+1)*16-1-:16];
                next_layer_0[9903-:16] = layer_0[9903-:16] + layer_input[9903-:16]*kernel_0[(39552+col+1)*16-1-:16];
                next_layer_0[9919-:16] = layer_0[9919-:16] + layer_input[9919-:16]*kernel_0[(39616+col+1)*16-1-:16];
                next_layer_0[9935-:16] = layer_0[9935-:16] + layer_input[9935-:16]*kernel_0[(39680+col+1)*16-1-:16];
                next_layer_0[9951-:16] = layer_0[9951-:16] + layer_input[9951-:16]*kernel_0[(39744+col+1)*16-1-:16];
                next_layer_0[9967-:16] = layer_0[9967-:16] + layer_input[9967-:16]*kernel_0[(39808+col+1)*16-1-:16];
                next_layer_0[9983-:16] = layer_0[9983-:16] + layer_input[9983-:16]*kernel_0[(39872+col+1)*16-1-:16];
                next_layer_0[9999-:16] = layer_0[9999-:16] + layer_input[9999-:16]*kernel_0[(39936+col+1)*16-1-:16];
                next_layer_0[10015-:16] = layer_0[10015-:16] + layer_input[10015-:16]*kernel_0[(40000+col+1)*16-1-:16];
                next_layer_0[10031-:16] = layer_0[10031-:16] + layer_input[10031-:16]*kernel_0[(40064+col+1)*16-1-:16];
                next_layer_0[10047-:16] = layer_0[10047-:16] + layer_input[10047-:16]*kernel_0[(40128+col+1)*16-1-:16];
                next_layer_0[10063-:16] = layer_0[10063-:16] + layer_input[10063-:16]*kernel_0[(40192+col+1)*16-1-:16];
                next_layer_0[10079-:16] = layer_0[10079-:16] + layer_input[10079-:16]*kernel_0[(40256+col+1)*16-1-:16];
                next_layer_0[10095-:16] = layer_0[10095-:16] + layer_input[10095-:16]*kernel_0[(40320+col+1)*16-1-:16];
                next_layer_0[10111-:16] = layer_0[10111-:16] + layer_input[10111-:16]*kernel_0[(40384+col+1)*16-1-:16];
                next_layer_0[10127-:16] = layer_0[10127-:16] + layer_input[10127-:16]*kernel_0[(40448+col+1)*16-1-:16];
                next_layer_0[10143-:16] = layer_0[10143-:16] + layer_input[10143-:16]*kernel_0[(40512+col+1)*16-1-:16];
                next_layer_0[10159-:16] = layer_0[10159-:16] + layer_input[10159-:16]*kernel_0[(40576+col+1)*16-1-:16];
                next_layer_0[10175-:16] = layer_0[10175-:16] + layer_input[10175-:16]*kernel_0[(40640+col+1)*16-1-:16];
                next_layer_0[10191-:16] = layer_0[10191-:16] + layer_input[10191-:16]*kernel_0[(40704+col+1)*16-1-:16];
                next_layer_0[10207-:16] = layer_0[10207-:16] + layer_input[10207-:16]*kernel_0[(40768+col+1)*16-1-:16];
                next_layer_0[10223-:16] = layer_0[10223-:16] + layer_input[10223-:16]*kernel_0[(40832+col+1)*16-1-:16];
                next_layer_0[10239-:16] = layer_0[10239-:16] + layer_input[10239-:16]*kernel_0[(40896+col+1)*16-1-:16];
                next_layer_0[10255-:16] = layer_0[10255-:16] + layer_input[10255-:16]*kernel_0[(40960+col+1)*16-1-:16];
                next_layer_0[10271-:16] = layer_0[10271-:16] + layer_input[10271-:16]*kernel_0[(41024+col+1)*16-1-:16];
                next_layer_0[10287-:16] = layer_0[10287-:16] + layer_input[10287-:16]*kernel_0[(41088+col+1)*16-1-:16];
                next_layer_0[10303-:16] = layer_0[10303-:16] + layer_input[10303-:16]*kernel_0[(41152+col+1)*16-1-:16];
                next_layer_0[10319-:16] = layer_0[10319-:16] + layer_input[10319-:16]*kernel_0[(41216+col+1)*16-1-:16];
                next_layer_0[10335-:16] = layer_0[10335-:16] + layer_input[10335-:16]*kernel_0[(41280+col+1)*16-1-:16];
                next_layer_0[10351-:16] = layer_0[10351-:16] + layer_input[10351-:16]*kernel_0[(41344+col+1)*16-1-:16];
                next_layer_0[10367-:16] = layer_0[10367-:16] + layer_input[10367-:16]*kernel_0[(41408+col+1)*16-1-:16];
                next_layer_0[10383-:16] = layer_0[10383-:16] + layer_input[10383-:16]*kernel_0[(41472+col+1)*16-1-:16];
                next_layer_0[10399-:16] = layer_0[10399-:16] + layer_input[10399-:16]*kernel_0[(41536+col+1)*16-1-:16];
                next_layer_0[10415-:16] = layer_0[10415-:16] + layer_input[10415-:16]*kernel_0[(41600+col+1)*16-1-:16];
                next_layer_0[10431-:16] = layer_0[10431-:16] + layer_input[10431-:16]*kernel_0[(41664+col+1)*16-1-:16];
                next_layer_0[10447-:16] = layer_0[10447-:16] + layer_input[10447-:16]*kernel_0[(41728+col+1)*16-1-:16];
                next_layer_0[10463-:16] = layer_0[10463-:16] + layer_input[10463-:16]*kernel_0[(41792+col+1)*16-1-:16];
                next_layer_0[10479-:16] = layer_0[10479-:16] + layer_input[10479-:16]*kernel_0[(41856+col+1)*16-1-:16];
                next_layer_0[10495-:16] = layer_0[10495-:16] + layer_input[10495-:16]*kernel_0[(41920+col+1)*16-1-:16];
                next_layer_0[10511-:16] = layer_0[10511-:16] + layer_input[10511-:16]*kernel_0[(41984+col+1)*16-1-:16];
                next_layer_0[10527-:16] = layer_0[10527-:16] + layer_input[10527-:16]*kernel_0[(42048+col+1)*16-1-:16];
                next_layer_0[10543-:16] = layer_0[10543-:16] + layer_input[10543-:16]*kernel_0[(42112+col+1)*16-1-:16];
                next_layer_0[10559-:16] = layer_0[10559-:16] + layer_input[10559-:16]*kernel_0[(42176+col+1)*16-1-:16];
                next_layer_0[10575-:16] = layer_0[10575-:16] + layer_input[10575-:16]*kernel_0[(42240+col+1)*16-1-:16];
                next_layer_0[10591-:16] = layer_0[10591-:16] + layer_input[10591-:16]*kernel_0[(42304+col+1)*16-1-:16];
                next_layer_0[10607-:16] = layer_0[10607-:16] + layer_input[10607-:16]*kernel_0[(42368+col+1)*16-1-:16];
                next_layer_0[10623-:16] = layer_0[10623-:16] + layer_input[10623-:16]*kernel_0[(42432+col+1)*16-1-:16];
                next_layer_0[10639-:16] = layer_0[10639-:16] + layer_input[10639-:16]*kernel_0[(42496+col+1)*16-1-:16];
                next_layer_0[10655-:16] = layer_0[10655-:16] + layer_input[10655-:16]*kernel_0[(42560+col+1)*16-1-:16];
                next_layer_0[10671-:16] = layer_0[10671-:16] + layer_input[10671-:16]*kernel_0[(42624+col+1)*16-1-:16];
                next_layer_0[10687-:16] = layer_0[10687-:16] + layer_input[10687-:16]*kernel_0[(42688+col+1)*16-1-:16];
                next_layer_0[10703-:16] = layer_0[10703-:16] + layer_input[10703-:16]*kernel_0[(42752+col+1)*16-1-:16];
                next_layer_0[10719-:16] = layer_0[10719-:16] + layer_input[10719-:16]*kernel_0[(42816+col+1)*16-1-:16];
                next_layer_0[10735-:16] = layer_0[10735-:16] + layer_input[10735-:16]*kernel_0[(42880+col+1)*16-1-:16];
                next_layer_0[10751-:16] = layer_0[10751-:16] + layer_input[10751-:16]*kernel_0[(42944+col+1)*16-1-:16];
                next_layer_0[10767-:16] = layer_0[10767-:16] + layer_input[10767-:16]*kernel_0[(43008+col+1)*16-1-:16];
                next_layer_0[10783-:16] = layer_0[10783-:16] + layer_input[10783-:16]*kernel_0[(43072+col+1)*16-1-:16];
                next_layer_0[10799-:16] = layer_0[10799-:16] + layer_input[10799-:16]*kernel_0[(43136+col+1)*16-1-:16];
                next_layer_0[10815-:16] = layer_0[10815-:16] + layer_input[10815-:16]*kernel_0[(43200+col+1)*16-1-:16];
                next_layer_0[10831-:16] = layer_0[10831-:16] + layer_input[10831-:16]*kernel_0[(43264+col+1)*16-1-:16];
                next_layer_0[10847-:16] = layer_0[10847-:16] + layer_input[10847-:16]*kernel_0[(43328+col+1)*16-1-:16];
                next_layer_0[10863-:16] = layer_0[10863-:16] + layer_input[10863-:16]*kernel_0[(43392+col+1)*16-1-:16];
                next_layer_0[10879-:16] = layer_0[10879-:16] + layer_input[10879-:16]*kernel_0[(43456+col+1)*16-1-:16];
                next_layer_0[10895-:16] = layer_0[10895-:16] + layer_input[10895-:16]*kernel_0[(43520+col+1)*16-1-:16];
                next_layer_0[10911-:16] = layer_0[10911-:16] + layer_input[10911-:16]*kernel_0[(43584+col+1)*16-1-:16];
                next_layer_0[10927-:16] = layer_0[10927-:16] + layer_input[10927-:16]*kernel_0[(43648+col+1)*16-1-:16];
                next_layer_0[10943-:16] = layer_0[10943-:16] + layer_input[10943-:16]*kernel_0[(43712+col+1)*16-1-:16];
                next_layer_0[10959-:16] = layer_0[10959-:16] + layer_input[10959-:16]*kernel_0[(43776+col+1)*16-1-:16];
                next_layer_0[10975-:16] = layer_0[10975-:16] + layer_input[10975-:16]*kernel_0[(43840+col+1)*16-1-:16];
                next_layer_0[10991-:16] = layer_0[10991-:16] + layer_input[10991-:16]*kernel_0[(43904+col+1)*16-1-:16];
                next_layer_0[11007-:16] = layer_0[11007-:16] + layer_input[11007-:16]*kernel_0[(43968+col+1)*16-1-:16];
                next_layer_0[11023-:16] = layer_0[11023-:16] + layer_input[11023-:16]*kernel_0[(44032+col+1)*16-1-:16];
                next_layer_0[11039-:16] = layer_0[11039-:16] + layer_input[11039-:16]*kernel_0[(44096+col+1)*16-1-:16];
                next_layer_0[11055-:16] = layer_0[11055-:16] + layer_input[11055-:16]*kernel_0[(44160+col+1)*16-1-:16];
                next_layer_0[11071-:16] = layer_0[11071-:16] + layer_input[11071-:16]*kernel_0[(44224+col+1)*16-1-:16];
                next_layer_0[11087-:16] = layer_0[11087-:16] + layer_input[11087-:16]*kernel_0[(44288+col+1)*16-1-:16];
                next_layer_0[11103-:16] = layer_0[11103-:16] + layer_input[11103-:16]*kernel_0[(44352+col+1)*16-1-:16];
                next_layer_0[11119-:16] = layer_0[11119-:16] + layer_input[11119-:16]*kernel_0[(44416+col+1)*16-1-:16];
                next_layer_0[11135-:16] = layer_0[11135-:16] + layer_input[11135-:16]*kernel_0[(44480+col+1)*16-1-:16];
                next_layer_0[11151-:16] = layer_0[11151-:16] + layer_input[11151-:16]*kernel_0[(44544+col+1)*16-1-:16];
                next_layer_0[11167-:16] = layer_0[11167-:16] + layer_input[11167-:16]*kernel_0[(44608+col+1)*16-1-:16];
                next_layer_0[11183-:16] = layer_0[11183-:16] + layer_input[11183-:16]*kernel_0[(44672+col+1)*16-1-:16];
                next_layer_0[11199-:16] = layer_0[11199-:16] + layer_input[11199-:16]*kernel_0[(44736+col+1)*16-1-:16];
                next_layer_0[11215-:16] = layer_0[11215-:16] + layer_input[11215-:16]*kernel_0[(44800+col+1)*16-1-:16];
                next_layer_0[11231-:16] = layer_0[11231-:16] + layer_input[11231-:16]*kernel_0[(44864+col+1)*16-1-:16];
                next_layer_0[11247-:16] = layer_0[11247-:16] + layer_input[11247-:16]*kernel_0[(44928+col+1)*16-1-:16];
                next_layer_0[11263-:16] = layer_0[11263-:16] + layer_input[11263-:16]*kernel_0[(44992+col+1)*16-1-:16];
                next_layer_0[11279-:16] = layer_0[11279-:16] + layer_input[11279-:16]*kernel_0[(45056+col+1)*16-1-:16];
                next_layer_0[11295-:16] = layer_0[11295-:16] + layer_input[11295-:16]*kernel_0[(45120+col+1)*16-1-:16];
                next_layer_0[11311-:16] = layer_0[11311-:16] + layer_input[11311-:16]*kernel_0[(45184+col+1)*16-1-:16];
                next_layer_0[11327-:16] = layer_0[11327-:16] + layer_input[11327-:16]*kernel_0[(45248+col+1)*16-1-:16];
                next_layer_0[11343-:16] = layer_0[11343-:16] + layer_input[11343-:16]*kernel_0[(45312+col+1)*16-1-:16];
                next_layer_0[11359-:16] = layer_0[11359-:16] + layer_input[11359-:16]*kernel_0[(45376+col+1)*16-1-:16];
                next_layer_0[11375-:16] = layer_0[11375-:16] + layer_input[11375-:16]*kernel_0[(45440+col+1)*16-1-:16];
                next_layer_0[11391-:16] = layer_0[11391-:16] + layer_input[11391-:16]*kernel_0[(45504+col+1)*16-1-:16];
                next_layer_0[11407-:16] = layer_0[11407-:16] + layer_input[11407-:16]*kernel_0[(45568+col+1)*16-1-:16];
                next_layer_0[11423-:16] = layer_0[11423-:16] + layer_input[11423-:16]*kernel_0[(45632+col+1)*16-1-:16];
                next_layer_0[11439-:16] = layer_0[11439-:16] + layer_input[11439-:16]*kernel_0[(45696+col+1)*16-1-:16];
                next_layer_0[11455-:16] = layer_0[11455-:16] + layer_input[11455-:16]*kernel_0[(45760+col+1)*16-1-:16];
                next_layer_0[11471-:16] = layer_0[11471-:16] + layer_input[11471-:16]*kernel_0[(45824+col+1)*16-1-:16];
                next_layer_0[11487-:16] = layer_0[11487-:16] + layer_input[11487-:16]*kernel_0[(45888+col+1)*16-1-:16];
                next_layer_0[11503-:16] = layer_0[11503-:16] + layer_input[11503-:16]*kernel_0[(45952+col+1)*16-1-:16];
                next_layer_0[11519-:16] = layer_0[11519-:16] + layer_input[11519-:16]*kernel_0[(46016+col+1)*16-1-:16];
                next_layer_0[11535-:16] = layer_0[11535-:16] + layer_input[11535-:16]*kernel_0[(46080+col+1)*16-1-:16];
                next_layer_0[11551-:16] = layer_0[11551-:16] + layer_input[11551-:16]*kernel_0[(46144+col+1)*16-1-:16];
                next_layer_0[11567-:16] = layer_0[11567-:16] + layer_input[11567-:16]*kernel_0[(46208+col+1)*16-1-:16];
                next_layer_0[11583-:16] = layer_0[11583-:16] + layer_input[11583-:16]*kernel_0[(46272+col+1)*16-1-:16];
                next_layer_0[11599-:16] = layer_0[11599-:16] + layer_input[11599-:16]*kernel_0[(46336+col+1)*16-1-:16];
                next_layer_0[11615-:16] = layer_0[11615-:16] + layer_input[11615-:16]*kernel_0[(46400+col+1)*16-1-:16];
                next_layer_0[11631-:16] = layer_0[11631-:16] + layer_input[11631-:16]*kernel_0[(46464+col+1)*16-1-:16];
                next_layer_0[11647-:16] = layer_0[11647-:16] + layer_input[11647-:16]*kernel_0[(46528+col+1)*16-1-:16];
                next_layer_0[11663-:16] = layer_0[11663-:16] + layer_input[11663-:16]*kernel_0[(46592+col+1)*16-1-:16];
                next_layer_0[11679-:16] = layer_0[11679-:16] + layer_input[11679-:16]*kernel_0[(46656+col+1)*16-1-:16];
                next_layer_0[11695-:16] = layer_0[11695-:16] + layer_input[11695-:16]*kernel_0[(46720+col+1)*16-1-:16];
                next_layer_0[11711-:16] = layer_0[11711-:16] + layer_input[11711-:16]*kernel_0[(46784+col+1)*16-1-:16];
                next_layer_0[11727-:16] = layer_0[11727-:16] + layer_input[11727-:16]*kernel_0[(46848+col+1)*16-1-:16];
                next_layer_0[11743-:16] = layer_0[11743-:16] + layer_input[11743-:16]*kernel_0[(46912+col+1)*16-1-:16];
                next_layer_0[11759-:16] = layer_0[11759-:16] + layer_input[11759-:16]*kernel_0[(46976+col+1)*16-1-:16];
                next_layer_0[11775-:16] = layer_0[11775-:16] + layer_input[11775-:16]*kernel_0[(47040+col+1)*16-1-:16];
                next_layer_0[11791-:16] = layer_0[11791-:16] + layer_input[11791-:16]*kernel_0[(47104+col+1)*16-1-:16];
                next_layer_0[11807-:16] = layer_0[11807-:16] + layer_input[11807-:16]*kernel_0[(47168+col+1)*16-1-:16];
                next_layer_0[11823-:16] = layer_0[11823-:16] + layer_input[11823-:16]*kernel_0[(47232+col+1)*16-1-:16];
                next_layer_0[11839-:16] = layer_0[11839-:16] + layer_input[11839-:16]*kernel_0[(47296+col+1)*16-1-:16];
                next_layer_0[11855-:16] = layer_0[11855-:16] + layer_input[11855-:16]*kernel_0[(47360+col+1)*16-1-:16];
                next_layer_0[11871-:16] = layer_0[11871-:16] + layer_input[11871-:16]*kernel_0[(47424+col+1)*16-1-:16];
                next_layer_0[11887-:16] = layer_0[11887-:16] + layer_input[11887-:16]*kernel_0[(47488+col+1)*16-1-:16];
                next_layer_0[11903-:16] = layer_0[11903-:16] + layer_input[11903-:16]*kernel_0[(47552+col+1)*16-1-:16];
                next_layer_0[11919-:16] = layer_0[11919-:16] + layer_input[11919-:16]*kernel_0[(47616+col+1)*16-1-:16];
                next_layer_0[11935-:16] = layer_0[11935-:16] + layer_input[11935-:16]*kernel_0[(47680+col+1)*16-1-:16];
                next_layer_0[11951-:16] = layer_0[11951-:16] + layer_input[11951-:16]*kernel_0[(47744+col+1)*16-1-:16];
                next_layer_0[11967-:16] = layer_0[11967-:16] + layer_input[11967-:16]*kernel_0[(47808+col+1)*16-1-:16];
                next_layer_0[11983-:16] = layer_0[11983-:16] + layer_input[11983-:16]*kernel_0[(47872+col+1)*16-1-:16];
                next_layer_0[11999-:16] = layer_0[11999-:16] + layer_input[11999-:16]*kernel_0[(47936+col+1)*16-1-:16];
                next_layer_0[12015-:16] = layer_0[12015-:16] + layer_input[12015-:16]*kernel_0[(48000+col+1)*16-1-:16];
                next_layer_0[12031-:16] = layer_0[12031-:16] + layer_input[12031-:16]*kernel_0[(48064+col+1)*16-1-:16];
                next_layer_0[12047-:16] = layer_0[12047-:16] + layer_input[12047-:16]*kernel_0[(48128+col+1)*16-1-:16];
                next_layer_0[12063-:16] = layer_0[12063-:16] + layer_input[12063-:16]*kernel_0[(48192+col+1)*16-1-:16];
                next_layer_0[12079-:16] = layer_0[12079-:16] + layer_input[12079-:16]*kernel_0[(48256+col+1)*16-1-:16];
                next_layer_0[12095-:16] = layer_0[12095-:16] + layer_input[12095-:16]*kernel_0[(48320+col+1)*16-1-:16];
                next_layer_0[12111-:16] = layer_0[12111-:16] + layer_input[12111-:16]*kernel_0[(48384+col+1)*16-1-:16];
                next_layer_0[12127-:16] = layer_0[12127-:16] + layer_input[12127-:16]*kernel_0[(48448+col+1)*16-1-:16];
                next_layer_0[12143-:16] = layer_0[12143-:16] + layer_input[12143-:16]*kernel_0[(48512+col+1)*16-1-:16];
                next_layer_0[12159-:16] = layer_0[12159-:16] + layer_input[12159-:16]*kernel_0[(48576+col+1)*16-1-:16];
                next_layer_0[12175-:16] = layer_0[12175-:16] + layer_input[12175-:16]*kernel_0[(48640+col+1)*16-1-:16];
                next_layer_0[12191-:16] = layer_0[12191-:16] + layer_input[12191-:16]*kernel_0[(48704+col+1)*16-1-:16];
                next_layer_0[12207-:16] = layer_0[12207-:16] + layer_input[12207-:16]*kernel_0[(48768+col+1)*16-1-:16];
                next_layer_0[12223-:16] = layer_0[12223-:16] + layer_input[12223-:16]*kernel_0[(48832+col+1)*16-1-:16];
                next_layer_0[12239-:16] = layer_0[12239-:16] + layer_input[12239-:16]*kernel_0[(48896+col+1)*16-1-:16];
                next_layer_0[12255-:16] = layer_0[12255-:16] + layer_input[12255-:16]*kernel_0[(48960+col+1)*16-1-:16];
                next_layer_0[12271-:16] = layer_0[12271-:16] + layer_input[12271-:16]*kernel_0[(49024+col+1)*16-1-:16];
                next_layer_0[12287-:16] = layer_0[12287-:16] + layer_input[12287-:16]*kernel_0[(49088+col+1)*16-1-:16];
                next_layer_0[12303-:16] = layer_0[12303-:16] + layer_input[12303-:16]*kernel_0[(49152+col+1)*16-1-:16];
                next_layer_0[12319-:16] = layer_0[12319-:16] + layer_input[12319-:16]*kernel_0[(49216+col+1)*16-1-:16];
                next_layer_0[12335-:16] = layer_0[12335-:16] + layer_input[12335-:16]*kernel_0[(49280+col+1)*16-1-:16];
                next_layer_0[12351-:16] = layer_0[12351-:16] + layer_input[12351-:16]*kernel_0[(49344+col+1)*16-1-:16];
                next_layer_0[12367-:16] = layer_0[12367-:16] + layer_input[12367-:16]*kernel_0[(49408+col+1)*16-1-:16];
                next_layer_0[12383-:16] = layer_0[12383-:16] + layer_input[12383-:16]*kernel_0[(49472+col+1)*16-1-:16];
                next_layer_0[12399-:16] = layer_0[12399-:16] + layer_input[12399-:16]*kernel_0[(49536+col+1)*16-1-:16];
                next_layer_0[12415-:16] = layer_0[12415-:16] + layer_input[12415-:16]*kernel_0[(49600+col+1)*16-1-:16];
                next_layer_0[12431-:16] = layer_0[12431-:16] + layer_input[12431-:16]*kernel_0[(49664+col+1)*16-1-:16];
                next_layer_0[12447-:16] = layer_0[12447-:16] + layer_input[12447-:16]*kernel_0[(49728+col+1)*16-1-:16];
                next_layer_0[12463-:16] = layer_0[12463-:16] + layer_input[12463-:16]*kernel_0[(49792+col+1)*16-1-:16];
                next_layer_0[12479-:16] = layer_0[12479-:16] + layer_input[12479-:16]*kernel_0[(49856+col+1)*16-1-:16];
                next_layer_0[12495-:16] = layer_0[12495-:16] + layer_input[12495-:16]*kernel_0[(49920+col+1)*16-1-:16];
                next_layer_0[12511-:16] = layer_0[12511-:16] + layer_input[12511-:16]*kernel_0[(49984+col+1)*16-1-:16];
                next_layer_0[12527-:16] = layer_0[12527-:16] + layer_input[12527-:16]*kernel_0[(50048+col+1)*16-1-:16];
                next_layer_0[12543-:16] = layer_0[12543-:16] + layer_input[12543-:16]*kernel_0[(50112+col+1)*16-1-:16];
            end
            SRELU: begin
                next_layer_0[15-:16] = (layer_0[15] ? -layer_0[15-:16] : layer_0[15-:16]);
                next_layer_0[31-:16] = (layer_0[31] ? -layer_0[31-:16] : layer_0[31-:16]);
                next_layer_0[47-:16] = (layer_0[47] ? -layer_0[47-:16] : layer_0[47-:16]);
                next_layer_0[63-:16] = (layer_0[63] ? -layer_0[63-:16] : layer_0[63-:16]);
                next_layer_0[79-:16] = (layer_0[79] ? -layer_0[79-:16] : layer_0[79-:16]);
                next_layer_0[95-:16] = (layer_0[95] ? -layer_0[95-:16] : layer_0[95-:16]);
                next_layer_0[111-:16] = (layer_0[111] ? -layer_0[111-:16] : layer_0[111-:16]);
                next_layer_0[127-:16] = (layer_0[127] ? -layer_0[127-:16] : layer_0[127-:16]);
                next_layer_0[143-:16] = (layer_0[143] ? -layer_0[143-:16] : layer_0[143-:16]);
                next_layer_0[159-:16] = (layer_0[159] ? -layer_0[159-:16] : layer_0[159-:16]);
                next_layer_0[175-:16] = (layer_0[175] ? -layer_0[175-:16] : layer_0[175-:16]);
                next_layer_0[191-:16] = (layer_0[191] ? -layer_0[191-:16] : layer_0[191-:16]);
                next_layer_0[207-:16] = (layer_0[207] ? -layer_0[207-:16] : layer_0[207-:16]);
                next_layer_0[223-:16] = (layer_0[223] ? -layer_0[223-:16] : layer_0[223-:16]);
                next_layer_0[239-:16] = (layer_0[239] ? -layer_0[239-:16] : layer_0[239-:16]);
                next_layer_0[255-:16] = (layer_0[255] ? -layer_0[255-:16] : layer_0[255-:16]);
                next_layer_0[271-:16] = (layer_0[271] ? -layer_0[271-:16] : layer_0[271-:16]);
                next_layer_0[287-:16] = (layer_0[287] ? -layer_0[287-:16] : layer_0[287-:16]);
                next_layer_0[303-:16] = (layer_0[303] ? -layer_0[303-:16] : layer_0[303-:16]);
                next_layer_0[319-:16] = (layer_0[319] ? -layer_0[319-:16] : layer_0[319-:16]);
                next_layer_0[335-:16] = (layer_0[335] ? -layer_0[335-:16] : layer_0[335-:16]);
                next_layer_0[351-:16] = (layer_0[351] ? -layer_0[351-:16] : layer_0[351-:16]);
                next_layer_0[367-:16] = (layer_0[367] ? -layer_0[367-:16] : layer_0[367-:16]);
                next_layer_0[383-:16] = (layer_0[383] ? -layer_0[383-:16] : layer_0[383-:16]);
                next_layer_0[399-:16] = (layer_0[399] ? -layer_0[399-:16] : layer_0[399-:16]);
                next_layer_0[415-:16] = (layer_0[415] ? -layer_0[415-:16] : layer_0[415-:16]);
                next_layer_0[431-:16] = (layer_0[431] ? -layer_0[431-:16] : layer_0[431-:16]);
                next_layer_0[447-:16] = (layer_0[447] ? -layer_0[447-:16] : layer_0[447-:16]);
                next_layer_0[463-:16] = (layer_0[463] ? -layer_0[463-:16] : layer_0[463-:16]);
                next_layer_0[479-:16] = (layer_0[479] ? -layer_0[479-:16] : layer_0[479-:16]);
                next_layer_0[495-:16] = (layer_0[495] ? -layer_0[495-:16] : layer_0[495-:16]);
                next_layer_0[511-:16] = (layer_0[511] ? -layer_0[511-:16] : layer_0[511-:16]);
                next_layer_0[527-:16] = (layer_0[527] ? -layer_0[527-:16] : layer_0[527-:16]);
                next_layer_0[543-:16] = (layer_0[543] ? -layer_0[543-:16] : layer_0[543-:16]);
                next_layer_0[559-:16] = (layer_0[559] ? -layer_0[559-:16] : layer_0[559-:16]);
                next_layer_0[575-:16] = (layer_0[575] ? -layer_0[575-:16] : layer_0[575-:16]);
                next_layer_0[591-:16] = (layer_0[591] ? -layer_0[591-:16] : layer_0[591-:16]);
                next_layer_0[607-:16] = (layer_0[607] ? -layer_0[607-:16] : layer_0[607-:16]);
                next_layer_0[623-:16] = (layer_0[623] ? -layer_0[623-:16] : layer_0[623-:16]);
                next_layer_0[639-:16] = (layer_0[639] ? -layer_0[639-:16] : layer_0[639-:16]);
                next_layer_0[655-:16] = (layer_0[655] ? -layer_0[655-:16] : layer_0[655-:16]);
                next_layer_0[671-:16] = (layer_0[671] ? -layer_0[671-:16] : layer_0[671-:16]);
                next_layer_0[687-:16] = (layer_0[687] ? -layer_0[687-:16] : layer_0[687-:16]);
                next_layer_0[703-:16] = (layer_0[703] ? -layer_0[703-:16] : layer_0[703-:16]);
                next_layer_0[719-:16] = (layer_0[719] ? -layer_0[719-:16] : layer_0[719-:16]);
                next_layer_0[735-:16] = (layer_0[735] ? -layer_0[735-:16] : layer_0[735-:16]);
                next_layer_0[751-:16] = (layer_0[751] ? -layer_0[751-:16] : layer_0[751-:16]);
                next_layer_0[767-:16] = (layer_0[767] ? -layer_0[767-:16] : layer_0[767-:16]);
                next_layer_0[783-:16] = (layer_0[783] ? -layer_0[783-:16] : layer_0[783-:16]);
                next_layer_0[799-:16] = (layer_0[799] ? -layer_0[799-:16] : layer_0[799-:16]);
                next_layer_0[815-:16] = (layer_0[815] ? -layer_0[815-:16] : layer_0[815-:16]);
                next_layer_0[831-:16] = (layer_0[831] ? -layer_0[831-:16] : layer_0[831-:16]);
                next_layer_0[847-:16] = (layer_0[847] ? -layer_0[847-:16] : layer_0[847-:16]);
                next_layer_0[863-:16] = (layer_0[863] ? -layer_0[863-:16] : layer_0[863-:16]);
                next_layer_0[879-:16] = (layer_0[879] ? -layer_0[879-:16] : layer_0[879-:16]);
                next_layer_0[895-:16] = (layer_0[895] ? -layer_0[895-:16] : layer_0[895-:16]);
                next_layer_0[911-:16] = (layer_0[911] ? -layer_0[911-:16] : layer_0[911-:16]);
                next_layer_0[927-:16] = (layer_0[927] ? -layer_0[927-:16] : layer_0[927-:16]);
                next_layer_0[943-:16] = (layer_0[943] ? -layer_0[943-:16] : layer_0[943-:16]);
                next_layer_0[959-:16] = (layer_0[959] ? -layer_0[959-:16] : layer_0[959-:16]);
                next_layer_0[975-:16] = (layer_0[975] ? -layer_0[975-:16] : layer_0[975-:16]);
                next_layer_0[991-:16] = (layer_0[991] ? -layer_0[991-:16] : layer_0[991-:16]);
                next_layer_0[1007-:16] = (layer_0[1007] ? -layer_0[1007-:16] : layer_0[1007-:16]);
                next_layer_0[1023-:16] = (layer_0[1023] ? -layer_0[1023-:16] : layer_0[1023-:16]);
                next_layer_0[1039-:16] = (layer_0[1039] ? -layer_0[1039-:16] : layer_0[1039-:16]);
                next_layer_0[1055-:16] = (layer_0[1055] ? -layer_0[1055-:16] : layer_0[1055-:16]);
                next_layer_0[1071-:16] = (layer_0[1071] ? -layer_0[1071-:16] : layer_0[1071-:16]);
                next_layer_0[1087-:16] = (layer_0[1087] ? -layer_0[1087-:16] : layer_0[1087-:16]);
                next_layer_0[1103-:16] = (layer_0[1103] ? -layer_0[1103-:16] : layer_0[1103-:16]);
                next_layer_0[1119-:16] = (layer_0[1119] ? -layer_0[1119-:16] : layer_0[1119-:16]);
                next_layer_0[1135-:16] = (layer_0[1135] ? -layer_0[1135-:16] : layer_0[1135-:16]);
                next_layer_0[1151-:16] = (layer_0[1151] ? -layer_0[1151-:16] : layer_0[1151-:16]);
                next_layer_0[1167-:16] = (layer_0[1167] ? -layer_0[1167-:16] : layer_0[1167-:16]);
                next_layer_0[1183-:16] = (layer_0[1183] ? -layer_0[1183-:16] : layer_0[1183-:16]);
                next_layer_0[1199-:16] = (layer_0[1199] ? -layer_0[1199-:16] : layer_0[1199-:16]);
                next_layer_0[1215-:16] = (layer_0[1215] ? -layer_0[1215-:16] : layer_0[1215-:16]);
                next_layer_0[1231-:16] = (layer_0[1231] ? -layer_0[1231-:16] : layer_0[1231-:16]);
                next_layer_0[1247-:16] = (layer_0[1247] ? -layer_0[1247-:16] : layer_0[1247-:16]);
                next_layer_0[1263-:16] = (layer_0[1263] ? -layer_0[1263-:16] : layer_0[1263-:16]);
                next_layer_0[1279-:16] = (layer_0[1279] ? -layer_0[1279-:16] : layer_0[1279-:16]);
                next_layer_0[1295-:16] = (layer_0[1295] ? -layer_0[1295-:16] : layer_0[1295-:16]);
                next_layer_0[1311-:16] = (layer_0[1311] ? -layer_0[1311-:16] : layer_0[1311-:16]);
                next_layer_0[1327-:16] = (layer_0[1327] ? -layer_0[1327-:16] : layer_0[1327-:16]);
                next_layer_0[1343-:16] = (layer_0[1343] ? -layer_0[1343-:16] : layer_0[1343-:16]);
                next_layer_0[1359-:16] = (layer_0[1359] ? -layer_0[1359-:16] : layer_0[1359-:16]);
                next_layer_0[1375-:16] = (layer_0[1375] ? -layer_0[1375-:16] : layer_0[1375-:16]);
                next_layer_0[1391-:16] = (layer_0[1391] ? -layer_0[1391-:16] : layer_0[1391-:16]);
                next_layer_0[1407-:16] = (layer_0[1407] ? -layer_0[1407-:16] : layer_0[1407-:16]);
                next_layer_0[1423-:16] = (layer_0[1423] ? -layer_0[1423-:16] : layer_0[1423-:16]);
                next_layer_0[1439-:16] = (layer_0[1439] ? -layer_0[1439-:16] : layer_0[1439-:16]);
                next_layer_0[1455-:16] = (layer_0[1455] ? -layer_0[1455-:16] : layer_0[1455-:16]);
                next_layer_0[1471-:16] = (layer_0[1471] ? -layer_0[1471-:16] : layer_0[1471-:16]);
                next_layer_0[1487-:16] = (layer_0[1487] ? -layer_0[1487-:16] : layer_0[1487-:16]);
                next_layer_0[1503-:16] = (layer_0[1503] ? -layer_0[1503-:16] : layer_0[1503-:16]);
                next_layer_0[1519-:16] = (layer_0[1519] ? -layer_0[1519-:16] : layer_0[1519-:16]);
                next_layer_0[1535-:16] = (layer_0[1535] ? -layer_0[1535-:16] : layer_0[1535-:16]);
                next_layer_0[1551-:16] = (layer_0[1551] ? -layer_0[1551-:16] : layer_0[1551-:16]);
                next_layer_0[1567-:16] = (layer_0[1567] ? -layer_0[1567-:16] : layer_0[1567-:16]);
                next_layer_0[1583-:16] = (layer_0[1583] ? -layer_0[1583-:16] : layer_0[1583-:16]);
                next_layer_0[1599-:16] = (layer_0[1599] ? -layer_0[1599-:16] : layer_0[1599-:16]);
                next_layer_0[1615-:16] = (layer_0[1615] ? -layer_0[1615-:16] : layer_0[1615-:16]);
                next_layer_0[1631-:16] = (layer_0[1631] ? -layer_0[1631-:16] : layer_0[1631-:16]);
                next_layer_0[1647-:16] = (layer_0[1647] ? -layer_0[1647-:16] : layer_0[1647-:16]);
                next_layer_0[1663-:16] = (layer_0[1663] ? -layer_0[1663-:16] : layer_0[1663-:16]);
                next_layer_0[1679-:16] = (layer_0[1679] ? -layer_0[1679-:16] : layer_0[1679-:16]);
                next_layer_0[1695-:16] = (layer_0[1695] ? -layer_0[1695-:16] : layer_0[1695-:16]);
                next_layer_0[1711-:16] = (layer_0[1711] ? -layer_0[1711-:16] : layer_0[1711-:16]);
                next_layer_0[1727-:16] = (layer_0[1727] ? -layer_0[1727-:16] : layer_0[1727-:16]);
                next_layer_0[1743-:16] = (layer_0[1743] ? -layer_0[1743-:16] : layer_0[1743-:16]);
                next_layer_0[1759-:16] = (layer_0[1759] ? -layer_0[1759-:16] : layer_0[1759-:16]);
                next_layer_0[1775-:16] = (layer_0[1775] ? -layer_0[1775-:16] : layer_0[1775-:16]);
                next_layer_0[1791-:16] = (layer_0[1791] ? -layer_0[1791-:16] : layer_0[1791-:16]);
                next_layer_0[1807-:16] = (layer_0[1807] ? -layer_0[1807-:16] : layer_0[1807-:16]);
                next_layer_0[1823-:16] = (layer_0[1823] ? -layer_0[1823-:16] : layer_0[1823-:16]);
                next_layer_0[1839-:16] = (layer_0[1839] ? -layer_0[1839-:16] : layer_0[1839-:16]);
                next_layer_0[1855-:16] = (layer_0[1855] ? -layer_0[1855-:16] : layer_0[1855-:16]);
                next_layer_0[1871-:16] = (layer_0[1871] ? -layer_0[1871-:16] : layer_0[1871-:16]);
                next_layer_0[1887-:16] = (layer_0[1887] ? -layer_0[1887-:16] : layer_0[1887-:16]);
                next_layer_0[1903-:16] = (layer_0[1903] ? -layer_0[1903-:16] : layer_0[1903-:16]);
                next_layer_0[1919-:16] = (layer_0[1919] ? -layer_0[1919-:16] : layer_0[1919-:16]);
                next_layer_0[1935-:16] = (layer_0[1935] ? -layer_0[1935-:16] : layer_0[1935-:16]);
                next_layer_0[1951-:16] = (layer_0[1951] ? -layer_0[1951-:16] : layer_0[1951-:16]);
                next_layer_0[1967-:16] = (layer_0[1967] ? -layer_0[1967-:16] : layer_0[1967-:16]);
                next_layer_0[1983-:16] = (layer_0[1983] ? -layer_0[1983-:16] : layer_0[1983-:16]);
                next_layer_0[1999-:16] = (layer_0[1999] ? -layer_0[1999-:16] : layer_0[1999-:16]);
                next_layer_0[2015-:16] = (layer_0[2015] ? -layer_0[2015-:16] : layer_0[2015-:16]);
                next_layer_0[2031-:16] = (layer_0[2031] ? -layer_0[2031-:16] : layer_0[2031-:16]);
                next_layer_0[2047-:16] = (layer_0[2047] ? -layer_0[2047-:16] : layer_0[2047-:16]);
                next_layer_0[2063-:16] = (layer_0[2063] ? -layer_0[2063-:16] : layer_0[2063-:16]);
                next_layer_0[2079-:16] = (layer_0[2079] ? -layer_0[2079-:16] : layer_0[2079-:16]);
                next_layer_0[2095-:16] = (layer_0[2095] ? -layer_0[2095-:16] : layer_0[2095-:16]);
                next_layer_0[2111-:16] = (layer_0[2111] ? -layer_0[2111-:16] : layer_0[2111-:16]);
                next_layer_0[2127-:16] = (layer_0[2127] ? -layer_0[2127-:16] : layer_0[2127-:16]);
                next_layer_0[2143-:16] = (layer_0[2143] ? -layer_0[2143-:16] : layer_0[2143-:16]);
                next_layer_0[2159-:16] = (layer_0[2159] ? -layer_0[2159-:16] : layer_0[2159-:16]);
                next_layer_0[2175-:16] = (layer_0[2175] ? -layer_0[2175-:16] : layer_0[2175-:16]);
                next_layer_0[2191-:16] = (layer_0[2191] ? -layer_0[2191-:16] : layer_0[2191-:16]);
                next_layer_0[2207-:16] = (layer_0[2207] ? -layer_0[2207-:16] : layer_0[2207-:16]);
                next_layer_0[2223-:16] = (layer_0[2223] ? -layer_0[2223-:16] : layer_0[2223-:16]);
                next_layer_0[2239-:16] = (layer_0[2239] ? -layer_0[2239-:16] : layer_0[2239-:16]);
                next_layer_0[2255-:16] = (layer_0[2255] ? -layer_0[2255-:16] : layer_0[2255-:16]);
                next_layer_0[2271-:16] = (layer_0[2271] ? -layer_0[2271-:16] : layer_0[2271-:16]);
                next_layer_0[2287-:16] = (layer_0[2287] ? -layer_0[2287-:16] : layer_0[2287-:16]);
                next_layer_0[2303-:16] = (layer_0[2303] ? -layer_0[2303-:16] : layer_0[2303-:16]);
                next_layer_0[2319-:16] = (layer_0[2319] ? -layer_0[2319-:16] : layer_0[2319-:16]);
                next_layer_0[2335-:16] = (layer_0[2335] ? -layer_0[2335-:16] : layer_0[2335-:16]);
                next_layer_0[2351-:16] = (layer_0[2351] ? -layer_0[2351-:16] : layer_0[2351-:16]);
                next_layer_0[2367-:16] = (layer_0[2367] ? -layer_0[2367-:16] : layer_0[2367-:16]);
                next_layer_0[2383-:16] = (layer_0[2383] ? -layer_0[2383-:16] : layer_0[2383-:16]);
                next_layer_0[2399-:16] = (layer_0[2399] ? -layer_0[2399-:16] : layer_0[2399-:16]);
                next_layer_0[2415-:16] = (layer_0[2415] ? -layer_0[2415-:16] : layer_0[2415-:16]);
                next_layer_0[2431-:16] = (layer_0[2431] ? -layer_0[2431-:16] : layer_0[2431-:16]);
                next_layer_0[2447-:16] = (layer_0[2447] ? -layer_0[2447-:16] : layer_0[2447-:16]);
                next_layer_0[2463-:16] = (layer_0[2463] ? -layer_0[2463-:16] : layer_0[2463-:16]);
                next_layer_0[2479-:16] = (layer_0[2479] ? -layer_0[2479-:16] : layer_0[2479-:16]);
                next_layer_0[2495-:16] = (layer_0[2495] ? -layer_0[2495-:16] : layer_0[2495-:16]);
                next_layer_0[2511-:16] = (layer_0[2511] ? -layer_0[2511-:16] : layer_0[2511-:16]);
                next_layer_0[2527-:16] = (layer_0[2527] ? -layer_0[2527-:16] : layer_0[2527-:16]);
                next_layer_0[2543-:16] = (layer_0[2543] ? -layer_0[2543-:16] : layer_0[2543-:16]);
                next_layer_0[2559-:16] = (layer_0[2559] ? -layer_0[2559-:16] : layer_0[2559-:16]);
                next_layer_0[2575-:16] = (layer_0[2575] ? -layer_0[2575-:16] : layer_0[2575-:16]);
                next_layer_0[2591-:16] = (layer_0[2591] ? -layer_0[2591-:16] : layer_0[2591-:16]);
                next_layer_0[2607-:16] = (layer_0[2607] ? -layer_0[2607-:16] : layer_0[2607-:16]);
                next_layer_0[2623-:16] = (layer_0[2623] ? -layer_0[2623-:16] : layer_0[2623-:16]);
                next_layer_0[2639-:16] = (layer_0[2639] ? -layer_0[2639-:16] : layer_0[2639-:16]);
                next_layer_0[2655-:16] = (layer_0[2655] ? -layer_0[2655-:16] : layer_0[2655-:16]);
                next_layer_0[2671-:16] = (layer_0[2671] ? -layer_0[2671-:16] : layer_0[2671-:16]);
                next_layer_0[2687-:16] = (layer_0[2687] ? -layer_0[2687-:16] : layer_0[2687-:16]);
                next_layer_0[2703-:16] = (layer_0[2703] ? -layer_0[2703-:16] : layer_0[2703-:16]);
                next_layer_0[2719-:16] = (layer_0[2719] ? -layer_0[2719-:16] : layer_0[2719-:16]);
                next_layer_0[2735-:16] = (layer_0[2735] ? -layer_0[2735-:16] : layer_0[2735-:16]);
                next_layer_0[2751-:16] = (layer_0[2751] ? -layer_0[2751-:16] : layer_0[2751-:16]);
                next_layer_0[2767-:16] = (layer_0[2767] ? -layer_0[2767-:16] : layer_0[2767-:16]);
                next_layer_0[2783-:16] = (layer_0[2783] ? -layer_0[2783-:16] : layer_0[2783-:16]);
                next_layer_0[2799-:16] = (layer_0[2799] ? -layer_0[2799-:16] : layer_0[2799-:16]);
                next_layer_0[2815-:16] = (layer_0[2815] ? -layer_0[2815-:16] : layer_0[2815-:16]);
                next_layer_0[2831-:16] = (layer_0[2831] ? -layer_0[2831-:16] : layer_0[2831-:16]);
                next_layer_0[2847-:16] = (layer_0[2847] ? -layer_0[2847-:16] : layer_0[2847-:16]);
                next_layer_0[2863-:16] = (layer_0[2863] ? -layer_0[2863-:16] : layer_0[2863-:16]);
                next_layer_0[2879-:16] = (layer_0[2879] ? -layer_0[2879-:16] : layer_0[2879-:16]);
                next_layer_0[2895-:16] = (layer_0[2895] ? -layer_0[2895-:16] : layer_0[2895-:16]);
                next_layer_0[2911-:16] = (layer_0[2911] ? -layer_0[2911-:16] : layer_0[2911-:16]);
                next_layer_0[2927-:16] = (layer_0[2927] ? -layer_0[2927-:16] : layer_0[2927-:16]);
                next_layer_0[2943-:16] = (layer_0[2943] ? -layer_0[2943-:16] : layer_0[2943-:16]);
                next_layer_0[2959-:16] = (layer_0[2959] ? -layer_0[2959-:16] : layer_0[2959-:16]);
                next_layer_0[2975-:16] = (layer_0[2975] ? -layer_0[2975-:16] : layer_0[2975-:16]);
                next_layer_0[2991-:16] = (layer_0[2991] ? -layer_0[2991-:16] : layer_0[2991-:16]);
                next_layer_0[3007-:16] = (layer_0[3007] ? -layer_0[3007-:16] : layer_0[3007-:16]);
                next_layer_0[3023-:16] = (layer_0[3023] ? -layer_0[3023-:16] : layer_0[3023-:16]);
                next_layer_0[3039-:16] = (layer_0[3039] ? -layer_0[3039-:16] : layer_0[3039-:16]);
                next_layer_0[3055-:16] = (layer_0[3055] ? -layer_0[3055-:16] : layer_0[3055-:16]);
                next_layer_0[3071-:16] = (layer_0[3071] ? -layer_0[3071-:16] : layer_0[3071-:16]);
                next_layer_0[3087-:16] = (layer_0[3087] ? -layer_0[3087-:16] : layer_0[3087-:16]);
                next_layer_0[3103-:16] = (layer_0[3103] ? -layer_0[3103-:16] : layer_0[3103-:16]);
                next_layer_0[3119-:16] = (layer_0[3119] ? -layer_0[3119-:16] : layer_0[3119-:16]);
                next_layer_0[3135-:16] = (layer_0[3135] ? -layer_0[3135-:16] : layer_0[3135-:16]);
                next_layer_0[3151-:16] = (layer_0[3151] ? -layer_0[3151-:16] : layer_0[3151-:16]);
                next_layer_0[3167-:16] = (layer_0[3167] ? -layer_0[3167-:16] : layer_0[3167-:16]);
                next_layer_0[3183-:16] = (layer_0[3183] ? -layer_0[3183-:16] : layer_0[3183-:16]);
                next_layer_0[3199-:16] = (layer_0[3199] ? -layer_0[3199-:16] : layer_0[3199-:16]);
                next_layer_0[3215-:16] = (layer_0[3215] ? -layer_0[3215-:16] : layer_0[3215-:16]);
                next_layer_0[3231-:16] = (layer_0[3231] ? -layer_0[3231-:16] : layer_0[3231-:16]);
                next_layer_0[3247-:16] = (layer_0[3247] ? -layer_0[3247-:16] : layer_0[3247-:16]);
                next_layer_0[3263-:16] = (layer_0[3263] ? -layer_0[3263-:16] : layer_0[3263-:16]);
                next_layer_0[3279-:16] = (layer_0[3279] ? -layer_0[3279-:16] : layer_0[3279-:16]);
                next_layer_0[3295-:16] = (layer_0[3295] ? -layer_0[3295-:16] : layer_0[3295-:16]);
                next_layer_0[3311-:16] = (layer_0[3311] ? -layer_0[3311-:16] : layer_0[3311-:16]);
                next_layer_0[3327-:16] = (layer_0[3327] ? -layer_0[3327-:16] : layer_0[3327-:16]);
                next_layer_0[3343-:16] = (layer_0[3343] ? -layer_0[3343-:16] : layer_0[3343-:16]);
                next_layer_0[3359-:16] = (layer_0[3359] ? -layer_0[3359-:16] : layer_0[3359-:16]);
                next_layer_0[3375-:16] = (layer_0[3375] ? -layer_0[3375-:16] : layer_0[3375-:16]);
                next_layer_0[3391-:16] = (layer_0[3391] ? -layer_0[3391-:16] : layer_0[3391-:16]);
                next_layer_0[3407-:16] = (layer_0[3407] ? -layer_0[3407-:16] : layer_0[3407-:16]);
                next_layer_0[3423-:16] = (layer_0[3423] ? -layer_0[3423-:16] : layer_0[3423-:16]);
                next_layer_0[3439-:16] = (layer_0[3439] ? -layer_0[3439-:16] : layer_0[3439-:16]);
                next_layer_0[3455-:16] = (layer_0[3455] ? -layer_0[3455-:16] : layer_0[3455-:16]);
                next_layer_0[3471-:16] = (layer_0[3471] ? -layer_0[3471-:16] : layer_0[3471-:16]);
                next_layer_0[3487-:16] = (layer_0[3487] ? -layer_0[3487-:16] : layer_0[3487-:16]);
                next_layer_0[3503-:16] = (layer_0[3503] ? -layer_0[3503-:16] : layer_0[3503-:16]);
                next_layer_0[3519-:16] = (layer_0[3519] ? -layer_0[3519-:16] : layer_0[3519-:16]);
                next_layer_0[3535-:16] = (layer_0[3535] ? -layer_0[3535-:16] : layer_0[3535-:16]);
                next_layer_0[3551-:16] = (layer_0[3551] ? -layer_0[3551-:16] : layer_0[3551-:16]);
                next_layer_0[3567-:16] = (layer_0[3567] ? -layer_0[3567-:16] : layer_0[3567-:16]);
                next_layer_0[3583-:16] = (layer_0[3583] ? -layer_0[3583-:16] : layer_0[3583-:16]);
                next_layer_0[3599-:16] = (layer_0[3599] ? -layer_0[3599-:16] : layer_0[3599-:16]);
                next_layer_0[3615-:16] = (layer_0[3615] ? -layer_0[3615-:16] : layer_0[3615-:16]);
                next_layer_0[3631-:16] = (layer_0[3631] ? -layer_0[3631-:16] : layer_0[3631-:16]);
                next_layer_0[3647-:16] = (layer_0[3647] ? -layer_0[3647-:16] : layer_0[3647-:16]);
                next_layer_0[3663-:16] = (layer_0[3663] ? -layer_0[3663-:16] : layer_0[3663-:16]);
                next_layer_0[3679-:16] = (layer_0[3679] ? -layer_0[3679-:16] : layer_0[3679-:16]);
                next_layer_0[3695-:16] = (layer_0[3695] ? -layer_0[3695-:16] : layer_0[3695-:16]);
                next_layer_0[3711-:16] = (layer_0[3711] ? -layer_0[3711-:16] : layer_0[3711-:16]);
                next_layer_0[3727-:16] = (layer_0[3727] ? -layer_0[3727-:16] : layer_0[3727-:16]);
                next_layer_0[3743-:16] = (layer_0[3743] ? -layer_0[3743-:16] : layer_0[3743-:16]);
                next_layer_0[3759-:16] = (layer_0[3759] ? -layer_0[3759-:16] : layer_0[3759-:16]);
                next_layer_0[3775-:16] = (layer_0[3775] ? -layer_0[3775-:16] : layer_0[3775-:16]);
                next_layer_0[3791-:16] = (layer_0[3791] ? -layer_0[3791-:16] : layer_0[3791-:16]);
                next_layer_0[3807-:16] = (layer_0[3807] ? -layer_0[3807-:16] : layer_0[3807-:16]);
                next_layer_0[3823-:16] = (layer_0[3823] ? -layer_0[3823-:16] : layer_0[3823-:16]);
                next_layer_0[3839-:16] = (layer_0[3839] ? -layer_0[3839-:16] : layer_0[3839-:16]);
                next_layer_0[3855-:16] = (layer_0[3855] ? -layer_0[3855-:16] : layer_0[3855-:16]);
                next_layer_0[3871-:16] = (layer_0[3871] ? -layer_0[3871-:16] : layer_0[3871-:16]);
                next_layer_0[3887-:16] = (layer_0[3887] ? -layer_0[3887-:16] : layer_0[3887-:16]);
                next_layer_0[3903-:16] = (layer_0[3903] ? -layer_0[3903-:16] : layer_0[3903-:16]);
                next_layer_0[3919-:16] = (layer_0[3919] ? -layer_0[3919-:16] : layer_0[3919-:16]);
                next_layer_0[3935-:16] = (layer_0[3935] ? -layer_0[3935-:16] : layer_0[3935-:16]);
                next_layer_0[3951-:16] = (layer_0[3951] ? -layer_0[3951-:16] : layer_0[3951-:16]);
                next_layer_0[3967-:16] = (layer_0[3967] ? -layer_0[3967-:16] : layer_0[3967-:16]);
                next_layer_0[3983-:16] = (layer_0[3983] ? -layer_0[3983-:16] : layer_0[3983-:16]);
                next_layer_0[3999-:16] = (layer_0[3999] ? -layer_0[3999-:16] : layer_0[3999-:16]);
                next_layer_0[4015-:16] = (layer_0[4015] ? -layer_0[4015-:16] : layer_0[4015-:16]);
                next_layer_0[4031-:16] = (layer_0[4031] ? -layer_0[4031-:16] : layer_0[4031-:16]);
                next_layer_0[4047-:16] = (layer_0[4047] ? -layer_0[4047-:16] : layer_0[4047-:16]);
                next_layer_0[4063-:16] = (layer_0[4063] ? -layer_0[4063-:16] : layer_0[4063-:16]);
                next_layer_0[4079-:16] = (layer_0[4079] ? -layer_0[4079-:16] : layer_0[4079-:16]);
                next_layer_0[4095-:16] = (layer_0[4095] ? -layer_0[4095-:16] : layer_0[4095-:16]);
                next_layer_0[4111-:16] = (layer_0[4111] ? -layer_0[4111-:16] : layer_0[4111-:16]);
                next_layer_0[4127-:16] = (layer_0[4127] ? -layer_0[4127-:16] : layer_0[4127-:16]);
                next_layer_0[4143-:16] = (layer_0[4143] ? -layer_0[4143-:16] : layer_0[4143-:16]);
                next_layer_0[4159-:16] = (layer_0[4159] ? -layer_0[4159-:16] : layer_0[4159-:16]);
                next_layer_0[4175-:16] = (layer_0[4175] ? -layer_0[4175-:16] : layer_0[4175-:16]);
                next_layer_0[4191-:16] = (layer_0[4191] ? -layer_0[4191-:16] : layer_0[4191-:16]);
                next_layer_0[4207-:16] = (layer_0[4207] ? -layer_0[4207-:16] : layer_0[4207-:16]);
                next_layer_0[4223-:16] = (layer_0[4223] ? -layer_0[4223-:16] : layer_0[4223-:16]);
                next_layer_0[4239-:16] = (layer_0[4239] ? -layer_0[4239-:16] : layer_0[4239-:16]);
                next_layer_0[4255-:16] = (layer_0[4255] ? -layer_0[4255-:16] : layer_0[4255-:16]);
                next_layer_0[4271-:16] = (layer_0[4271] ? -layer_0[4271-:16] : layer_0[4271-:16]);
                next_layer_0[4287-:16] = (layer_0[4287] ? -layer_0[4287-:16] : layer_0[4287-:16]);
                next_layer_0[4303-:16] = (layer_0[4303] ? -layer_0[4303-:16] : layer_0[4303-:16]);
                next_layer_0[4319-:16] = (layer_0[4319] ? -layer_0[4319-:16] : layer_0[4319-:16]);
                next_layer_0[4335-:16] = (layer_0[4335] ? -layer_0[4335-:16] : layer_0[4335-:16]);
                next_layer_0[4351-:16] = (layer_0[4351] ? -layer_0[4351-:16] : layer_0[4351-:16]);
                next_layer_0[4367-:16] = (layer_0[4367] ? -layer_0[4367-:16] : layer_0[4367-:16]);
                next_layer_0[4383-:16] = (layer_0[4383] ? -layer_0[4383-:16] : layer_0[4383-:16]);
                next_layer_0[4399-:16] = (layer_0[4399] ? -layer_0[4399-:16] : layer_0[4399-:16]);
                next_layer_0[4415-:16] = (layer_0[4415] ? -layer_0[4415-:16] : layer_0[4415-:16]);
                next_layer_0[4431-:16] = (layer_0[4431] ? -layer_0[4431-:16] : layer_0[4431-:16]);
                next_layer_0[4447-:16] = (layer_0[4447] ? -layer_0[4447-:16] : layer_0[4447-:16]);
                next_layer_0[4463-:16] = (layer_0[4463] ? -layer_0[4463-:16] : layer_0[4463-:16]);
                next_layer_0[4479-:16] = (layer_0[4479] ? -layer_0[4479-:16] : layer_0[4479-:16]);
                next_layer_0[4495-:16] = (layer_0[4495] ? -layer_0[4495-:16] : layer_0[4495-:16]);
                next_layer_0[4511-:16] = (layer_0[4511] ? -layer_0[4511-:16] : layer_0[4511-:16]);
                next_layer_0[4527-:16] = (layer_0[4527] ? -layer_0[4527-:16] : layer_0[4527-:16]);
                next_layer_0[4543-:16] = (layer_0[4543] ? -layer_0[4543-:16] : layer_0[4543-:16]);
                next_layer_0[4559-:16] = (layer_0[4559] ? -layer_0[4559-:16] : layer_0[4559-:16]);
                next_layer_0[4575-:16] = (layer_0[4575] ? -layer_0[4575-:16] : layer_0[4575-:16]);
                next_layer_0[4591-:16] = (layer_0[4591] ? -layer_0[4591-:16] : layer_0[4591-:16]);
                next_layer_0[4607-:16] = (layer_0[4607] ? -layer_0[4607-:16] : layer_0[4607-:16]);
                next_layer_0[4623-:16] = (layer_0[4623] ? -layer_0[4623-:16] : layer_0[4623-:16]);
                next_layer_0[4639-:16] = (layer_0[4639] ? -layer_0[4639-:16] : layer_0[4639-:16]);
                next_layer_0[4655-:16] = (layer_0[4655] ? -layer_0[4655-:16] : layer_0[4655-:16]);
                next_layer_0[4671-:16] = (layer_0[4671] ? -layer_0[4671-:16] : layer_0[4671-:16]);
                next_layer_0[4687-:16] = (layer_0[4687] ? -layer_0[4687-:16] : layer_0[4687-:16]);
                next_layer_0[4703-:16] = (layer_0[4703] ? -layer_0[4703-:16] : layer_0[4703-:16]);
                next_layer_0[4719-:16] = (layer_0[4719] ? -layer_0[4719-:16] : layer_0[4719-:16]);
                next_layer_0[4735-:16] = (layer_0[4735] ? -layer_0[4735-:16] : layer_0[4735-:16]);
                next_layer_0[4751-:16] = (layer_0[4751] ? -layer_0[4751-:16] : layer_0[4751-:16]);
                next_layer_0[4767-:16] = (layer_0[4767] ? -layer_0[4767-:16] : layer_0[4767-:16]);
                next_layer_0[4783-:16] = (layer_0[4783] ? -layer_0[4783-:16] : layer_0[4783-:16]);
                next_layer_0[4799-:16] = (layer_0[4799] ? -layer_0[4799-:16] : layer_0[4799-:16]);
                next_layer_0[4815-:16] = (layer_0[4815] ? -layer_0[4815-:16] : layer_0[4815-:16]);
                next_layer_0[4831-:16] = (layer_0[4831] ? -layer_0[4831-:16] : layer_0[4831-:16]);
                next_layer_0[4847-:16] = (layer_0[4847] ? -layer_0[4847-:16] : layer_0[4847-:16]);
                next_layer_0[4863-:16] = (layer_0[4863] ? -layer_0[4863-:16] : layer_0[4863-:16]);
                next_layer_0[4879-:16] = (layer_0[4879] ? -layer_0[4879-:16] : layer_0[4879-:16]);
                next_layer_0[4895-:16] = (layer_0[4895] ? -layer_0[4895-:16] : layer_0[4895-:16]);
                next_layer_0[4911-:16] = (layer_0[4911] ? -layer_0[4911-:16] : layer_0[4911-:16]);
                next_layer_0[4927-:16] = (layer_0[4927] ? -layer_0[4927-:16] : layer_0[4927-:16]);
                next_layer_0[4943-:16] = (layer_0[4943] ? -layer_0[4943-:16] : layer_0[4943-:16]);
                next_layer_0[4959-:16] = (layer_0[4959] ? -layer_0[4959-:16] : layer_0[4959-:16]);
                next_layer_0[4975-:16] = (layer_0[4975] ? -layer_0[4975-:16] : layer_0[4975-:16]);
                next_layer_0[4991-:16] = (layer_0[4991] ? -layer_0[4991-:16] : layer_0[4991-:16]);
                next_layer_0[5007-:16] = (layer_0[5007] ? -layer_0[5007-:16] : layer_0[5007-:16]);
                next_layer_0[5023-:16] = (layer_0[5023] ? -layer_0[5023-:16] : layer_0[5023-:16]);
                next_layer_0[5039-:16] = (layer_0[5039] ? -layer_0[5039-:16] : layer_0[5039-:16]);
                next_layer_0[5055-:16] = (layer_0[5055] ? -layer_0[5055-:16] : layer_0[5055-:16]);
                next_layer_0[5071-:16] = (layer_0[5071] ? -layer_0[5071-:16] : layer_0[5071-:16]);
                next_layer_0[5087-:16] = (layer_0[5087] ? -layer_0[5087-:16] : layer_0[5087-:16]);
                next_layer_0[5103-:16] = (layer_0[5103] ? -layer_0[5103-:16] : layer_0[5103-:16]);
                next_layer_0[5119-:16] = (layer_0[5119] ? -layer_0[5119-:16] : layer_0[5119-:16]);
                next_layer_0[5135-:16] = (layer_0[5135] ? -layer_0[5135-:16] : layer_0[5135-:16]);
                next_layer_0[5151-:16] = (layer_0[5151] ? -layer_0[5151-:16] : layer_0[5151-:16]);
                next_layer_0[5167-:16] = (layer_0[5167] ? -layer_0[5167-:16] : layer_0[5167-:16]);
                next_layer_0[5183-:16] = (layer_0[5183] ? -layer_0[5183-:16] : layer_0[5183-:16]);
                next_layer_0[5199-:16] = (layer_0[5199] ? -layer_0[5199-:16] : layer_0[5199-:16]);
                next_layer_0[5215-:16] = (layer_0[5215] ? -layer_0[5215-:16] : layer_0[5215-:16]);
                next_layer_0[5231-:16] = (layer_0[5231] ? -layer_0[5231-:16] : layer_0[5231-:16]);
                next_layer_0[5247-:16] = (layer_0[5247] ? -layer_0[5247-:16] : layer_0[5247-:16]);
                next_layer_0[5263-:16] = (layer_0[5263] ? -layer_0[5263-:16] : layer_0[5263-:16]);
                next_layer_0[5279-:16] = (layer_0[5279] ? -layer_0[5279-:16] : layer_0[5279-:16]);
                next_layer_0[5295-:16] = (layer_0[5295] ? -layer_0[5295-:16] : layer_0[5295-:16]);
                next_layer_0[5311-:16] = (layer_0[5311] ? -layer_0[5311-:16] : layer_0[5311-:16]);
                next_layer_0[5327-:16] = (layer_0[5327] ? -layer_0[5327-:16] : layer_0[5327-:16]);
                next_layer_0[5343-:16] = (layer_0[5343] ? -layer_0[5343-:16] : layer_0[5343-:16]);
                next_layer_0[5359-:16] = (layer_0[5359] ? -layer_0[5359-:16] : layer_0[5359-:16]);
                next_layer_0[5375-:16] = (layer_0[5375] ? -layer_0[5375-:16] : layer_0[5375-:16]);
                next_layer_0[5391-:16] = (layer_0[5391] ? -layer_0[5391-:16] : layer_0[5391-:16]);
                next_layer_0[5407-:16] = (layer_0[5407] ? -layer_0[5407-:16] : layer_0[5407-:16]);
                next_layer_0[5423-:16] = (layer_0[5423] ? -layer_0[5423-:16] : layer_0[5423-:16]);
                next_layer_0[5439-:16] = (layer_0[5439] ? -layer_0[5439-:16] : layer_0[5439-:16]);
                next_layer_0[5455-:16] = (layer_0[5455] ? -layer_0[5455-:16] : layer_0[5455-:16]);
                next_layer_0[5471-:16] = (layer_0[5471] ? -layer_0[5471-:16] : layer_0[5471-:16]);
                next_layer_0[5487-:16] = (layer_0[5487] ? -layer_0[5487-:16] : layer_0[5487-:16]);
                next_layer_0[5503-:16] = (layer_0[5503] ? -layer_0[5503-:16] : layer_0[5503-:16]);
                next_layer_0[5519-:16] = (layer_0[5519] ? -layer_0[5519-:16] : layer_0[5519-:16]);
                next_layer_0[5535-:16] = (layer_0[5535] ? -layer_0[5535-:16] : layer_0[5535-:16]);
                next_layer_0[5551-:16] = (layer_0[5551] ? -layer_0[5551-:16] : layer_0[5551-:16]);
                next_layer_0[5567-:16] = (layer_0[5567] ? -layer_0[5567-:16] : layer_0[5567-:16]);
                next_layer_0[5583-:16] = (layer_0[5583] ? -layer_0[5583-:16] : layer_0[5583-:16]);
                next_layer_0[5599-:16] = (layer_0[5599] ? -layer_0[5599-:16] : layer_0[5599-:16]);
                next_layer_0[5615-:16] = (layer_0[5615] ? -layer_0[5615-:16] : layer_0[5615-:16]);
                next_layer_0[5631-:16] = (layer_0[5631] ? -layer_0[5631-:16] : layer_0[5631-:16]);
                next_layer_0[5647-:16] = (layer_0[5647] ? -layer_0[5647-:16] : layer_0[5647-:16]);
                next_layer_0[5663-:16] = (layer_0[5663] ? -layer_0[5663-:16] : layer_0[5663-:16]);
                next_layer_0[5679-:16] = (layer_0[5679] ? -layer_0[5679-:16] : layer_0[5679-:16]);
                next_layer_0[5695-:16] = (layer_0[5695] ? -layer_0[5695-:16] : layer_0[5695-:16]);
                next_layer_0[5711-:16] = (layer_0[5711] ? -layer_0[5711-:16] : layer_0[5711-:16]);
                next_layer_0[5727-:16] = (layer_0[5727] ? -layer_0[5727-:16] : layer_0[5727-:16]);
                next_layer_0[5743-:16] = (layer_0[5743] ? -layer_0[5743-:16] : layer_0[5743-:16]);
                next_layer_0[5759-:16] = (layer_0[5759] ? -layer_0[5759-:16] : layer_0[5759-:16]);
                next_layer_0[5775-:16] = (layer_0[5775] ? -layer_0[5775-:16] : layer_0[5775-:16]);
                next_layer_0[5791-:16] = (layer_0[5791] ? -layer_0[5791-:16] : layer_0[5791-:16]);
                next_layer_0[5807-:16] = (layer_0[5807] ? -layer_0[5807-:16] : layer_0[5807-:16]);
                next_layer_0[5823-:16] = (layer_0[5823] ? -layer_0[5823-:16] : layer_0[5823-:16]);
                next_layer_0[5839-:16] = (layer_0[5839] ? -layer_0[5839-:16] : layer_0[5839-:16]);
                next_layer_0[5855-:16] = (layer_0[5855] ? -layer_0[5855-:16] : layer_0[5855-:16]);
                next_layer_0[5871-:16] = (layer_0[5871] ? -layer_0[5871-:16] : layer_0[5871-:16]);
                next_layer_0[5887-:16] = (layer_0[5887] ? -layer_0[5887-:16] : layer_0[5887-:16]);
                next_layer_0[5903-:16] = (layer_0[5903] ? -layer_0[5903-:16] : layer_0[5903-:16]);
                next_layer_0[5919-:16] = (layer_0[5919] ? -layer_0[5919-:16] : layer_0[5919-:16]);
                next_layer_0[5935-:16] = (layer_0[5935] ? -layer_0[5935-:16] : layer_0[5935-:16]);
                next_layer_0[5951-:16] = (layer_0[5951] ? -layer_0[5951-:16] : layer_0[5951-:16]);
                next_layer_0[5967-:16] = (layer_0[5967] ? -layer_0[5967-:16] : layer_0[5967-:16]);
                next_layer_0[5983-:16] = (layer_0[5983] ? -layer_0[5983-:16] : layer_0[5983-:16]);
                next_layer_0[5999-:16] = (layer_0[5999] ? -layer_0[5999-:16] : layer_0[5999-:16]);
                next_layer_0[6015-:16] = (layer_0[6015] ? -layer_0[6015-:16] : layer_0[6015-:16]);
                next_layer_0[6031-:16] = (layer_0[6031] ? -layer_0[6031-:16] : layer_0[6031-:16]);
                next_layer_0[6047-:16] = (layer_0[6047] ? -layer_0[6047-:16] : layer_0[6047-:16]);
                next_layer_0[6063-:16] = (layer_0[6063] ? -layer_0[6063-:16] : layer_0[6063-:16]);
                next_layer_0[6079-:16] = (layer_0[6079] ? -layer_0[6079-:16] : layer_0[6079-:16]);
                next_layer_0[6095-:16] = (layer_0[6095] ? -layer_0[6095-:16] : layer_0[6095-:16]);
                next_layer_0[6111-:16] = (layer_0[6111] ? -layer_0[6111-:16] : layer_0[6111-:16]);
                next_layer_0[6127-:16] = (layer_0[6127] ? -layer_0[6127-:16] : layer_0[6127-:16]);
                next_layer_0[6143-:16] = (layer_0[6143] ? -layer_0[6143-:16] : layer_0[6143-:16]);
                next_layer_0[6159-:16] = (layer_0[6159] ? -layer_0[6159-:16] : layer_0[6159-:16]);
                next_layer_0[6175-:16] = (layer_0[6175] ? -layer_0[6175-:16] : layer_0[6175-:16]);
                next_layer_0[6191-:16] = (layer_0[6191] ? -layer_0[6191-:16] : layer_0[6191-:16]);
                next_layer_0[6207-:16] = (layer_0[6207] ? -layer_0[6207-:16] : layer_0[6207-:16]);
                next_layer_0[6223-:16] = (layer_0[6223] ? -layer_0[6223-:16] : layer_0[6223-:16]);
                next_layer_0[6239-:16] = (layer_0[6239] ? -layer_0[6239-:16] : layer_0[6239-:16]);
                next_layer_0[6255-:16] = (layer_0[6255] ? -layer_0[6255-:16] : layer_0[6255-:16]);
                next_layer_0[6271-:16] = (layer_0[6271] ? -layer_0[6271-:16] : layer_0[6271-:16]);
                next_layer_0[6287-:16] = (layer_0[6287] ? -layer_0[6287-:16] : layer_0[6287-:16]);
                next_layer_0[6303-:16] = (layer_0[6303] ? -layer_0[6303-:16] : layer_0[6303-:16]);
                next_layer_0[6319-:16] = (layer_0[6319] ? -layer_0[6319-:16] : layer_0[6319-:16]);
                next_layer_0[6335-:16] = (layer_0[6335] ? -layer_0[6335-:16] : layer_0[6335-:16]);
                next_layer_0[6351-:16] = (layer_0[6351] ? -layer_0[6351-:16] : layer_0[6351-:16]);
                next_layer_0[6367-:16] = (layer_0[6367] ? -layer_0[6367-:16] : layer_0[6367-:16]);
                next_layer_0[6383-:16] = (layer_0[6383] ? -layer_0[6383-:16] : layer_0[6383-:16]);
                next_layer_0[6399-:16] = (layer_0[6399] ? -layer_0[6399-:16] : layer_0[6399-:16]);
                next_layer_0[6415-:16] = (layer_0[6415] ? -layer_0[6415-:16] : layer_0[6415-:16]);
                next_layer_0[6431-:16] = (layer_0[6431] ? -layer_0[6431-:16] : layer_0[6431-:16]);
                next_layer_0[6447-:16] = (layer_0[6447] ? -layer_0[6447-:16] : layer_0[6447-:16]);
                next_layer_0[6463-:16] = (layer_0[6463] ? -layer_0[6463-:16] : layer_0[6463-:16]);
                next_layer_0[6479-:16] = (layer_0[6479] ? -layer_0[6479-:16] : layer_0[6479-:16]);
                next_layer_0[6495-:16] = (layer_0[6495] ? -layer_0[6495-:16] : layer_0[6495-:16]);
                next_layer_0[6511-:16] = (layer_0[6511] ? -layer_0[6511-:16] : layer_0[6511-:16]);
                next_layer_0[6527-:16] = (layer_0[6527] ? -layer_0[6527-:16] : layer_0[6527-:16]);
                next_layer_0[6543-:16] = (layer_0[6543] ? -layer_0[6543-:16] : layer_0[6543-:16]);
                next_layer_0[6559-:16] = (layer_0[6559] ? -layer_0[6559-:16] : layer_0[6559-:16]);
                next_layer_0[6575-:16] = (layer_0[6575] ? -layer_0[6575-:16] : layer_0[6575-:16]);
                next_layer_0[6591-:16] = (layer_0[6591] ? -layer_0[6591-:16] : layer_0[6591-:16]);
                next_layer_0[6607-:16] = (layer_0[6607] ? -layer_0[6607-:16] : layer_0[6607-:16]);
                next_layer_0[6623-:16] = (layer_0[6623] ? -layer_0[6623-:16] : layer_0[6623-:16]);
                next_layer_0[6639-:16] = (layer_0[6639] ? -layer_0[6639-:16] : layer_0[6639-:16]);
                next_layer_0[6655-:16] = (layer_0[6655] ? -layer_0[6655-:16] : layer_0[6655-:16]);
                next_layer_0[6671-:16] = (layer_0[6671] ? -layer_0[6671-:16] : layer_0[6671-:16]);
                next_layer_0[6687-:16] = (layer_0[6687] ? -layer_0[6687-:16] : layer_0[6687-:16]);
                next_layer_0[6703-:16] = (layer_0[6703] ? -layer_0[6703-:16] : layer_0[6703-:16]);
                next_layer_0[6719-:16] = (layer_0[6719] ? -layer_0[6719-:16] : layer_0[6719-:16]);
                next_layer_0[6735-:16] = (layer_0[6735] ? -layer_0[6735-:16] : layer_0[6735-:16]);
                next_layer_0[6751-:16] = (layer_0[6751] ? -layer_0[6751-:16] : layer_0[6751-:16]);
                next_layer_0[6767-:16] = (layer_0[6767] ? -layer_0[6767-:16] : layer_0[6767-:16]);
                next_layer_0[6783-:16] = (layer_0[6783] ? -layer_0[6783-:16] : layer_0[6783-:16]);
                next_layer_0[6799-:16] = (layer_0[6799] ? -layer_0[6799-:16] : layer_0[6799-:16]);
                next_layer_0[6815-:16] = (layer_0[6815] ? -layer_0[6815-:16] : layer_0[6815-:16]);
                next_layer_0[6831-:16] = (layer_0[6831] ? -layer_0[6831-:16] : layer_0[6831-:16]);
                next_layer_0[6847-:16] = (layer_0[6847] ? -layer_0[6847-:16] : layer_0[6847-:16]);
                next_layer_0[6863-:16] = (layer_0[6863] ? -layer_0[6863-:16] : layer_0[6863-:16]);
                next_layer_0[6879-:16] = (layer_0[6879] ? -layer_0[6879-:16] : layer_0[6879-:16]);
                next_layer_0[6895-:16] = (layer_0[6895] ? -layer_0[6895-:16] : layer_0[6895-:16]);
                next_layer_0[6911-:16] = (layer_0[6911] ? -layer_0[6911-:16] : layer_0[6911-:16]);
                next_layer_0[6927-:16] = (layer_0[6927] ? -layer_0[6927-:16] : layer_0[6927-:16]);
                next_layer_0[6943-:16] = (layer_0[6943] ? -layer_0[6943-:16] : layer_0[6943-:16]);
                next_layer_0[6959-:16] = (layer_0[6959] ? -layer_0[6959-:16] : layer_0[6959-:16]);
                next_layer_0[6975-:16] = (layer_0[6975] ? -layer_0[6975-:16] : layer_0[6975-:16]);
                next_layer_0[6991-:16] = (layer_0[6991] ? -layer_0[6991-:16] : layer_0[6991-:16]);
                next_layer_0[7007-:16] = (layer_0[7007] ? -layer_0[7007-:16] : layer_0[7007-:16]);
                next_layer_0[7023-:16] = (layer_0[7023] ? -layer_0[7023-:16] : layer_0[7023-:16]);
                next_layer_0[7039-:16] = (layer_0[7039] ? -layer_0[7039-:16] : layer_0[7039-:16]);
                next_layer_0[7055-:16] = (layer_0[7055] ? -layer_0[7055-:16] : layer_0[7055-:16]);
                next_layer_0[7071-:16] = (layer_0[7071] ? -layer_0[7071-:16] : layer_0[7071-:16]);
                next_layer_0[7087-:16] = (layer_0[7087] ? -layer_0[7087-:16] : layer_0[7087-:16]);
                next_layer_0[7103-:16] = (layer_0[7103] ? -layer_0[7103-:16] : layer_0[7103-:16]);
                next_layer_0[7119-:16] = (layer_0[7119] ? -layer_0[7119-:16] : layer_0[7119-:16]);
                next_layer_0[7135-:16] = (layer_0[7135] ? -layer_0[7135-:16] : layer_0[7135-:16]);
                next_layer_0[7151-:16] = (layer_0[7151] ? -layer_0[7151-:16] : layer_0[7151-:16]);
                next_layer_0[7167-:16] = (layer_0[7167] ? -layer_0[7167-:16] : layer_0[7167-:16]);
                next_layer_0[7183-:16] = (layer_0[7183] ? -layer_0[7183-:16] : layer_0[7183-:16]);
                next_layer_0[7199-:16] = (layer_0[7199] ? -layer_0[7199-:16] : layer_0[7199-:16]);
                next_layer_0[7215-:16] = (layer_0[7215] ? -layer_0[7215-:16] : layer_0[7215-:16]);
                next_layer_0[7231-:16] = (layer_0[7231] ? -layer_0[7231-:16] : layer_0[7231-:16]);
                next_layer_0[7247-:16] = (layer_0[7247] ? -layer_0[7247-:16] : layer_0[7247-:16]);
                next_layer_0[7263-:16] = (layer_0[7263] ? -layer_0[7263-:16] : layer_0[7263-:16]);
                next_layer_0[7279-:16] = (layer_0[7279] ? -layer_0[7279-:16] : layer_0[7279-:16]);
                next_layer_0[7295-:16] = (layer_0[7295] ? -layer_0[7295-:16] : layer_0[7295-:16]);
                next_layer_0[7311-:16] = (layer_0[7311] ? -layer_0[7311-:16] : layer_0[7311-:16]);
                next_layer_0[7327-:16] = (layer_0[7327] ? -layer_0[7327-:16] : layer_0[7327-:16]);
                next_layer_0[7343-:16] = (layer_0[7343] ? -layer_0[7343-:16] : layer_0[7343-:16]);
                next_layer_0[7359-:16] = (layer_0[7359] ? -layer_0[7359-:16] : layer_0[7359-:16]);
                next_layer_0[7375-:16] = (layer_0[7375] ? -layer_0[7375-:16] : layer_0[7375-:16]);
                next_layer_0[7391-:16] = (layer_0[7391] ? -layer_0[7391-:16] : layer_0[7391-:16]);
                next_layer_0[7407-:16] = (layer_0[7407] ? -layer_0[7407-:16] : layer_0[7407-:16]);
                next_layer_0[7423-:16] = (layer_0[7423] ? -layer_0[7423-:16] : layer_0[7423-:16]);
                next_layer_0[7439-:16] = (layer_0[7439] ? -layer_0[7439-:16] : layer_0[7439-:16]);
                next_layer_0[7455-:16] = (layer_0[7455] ? -layer_0[7455-:16] : layer_0[7455-:16]);
                next_layer_0[7471-:16] = (layer_0[7471] ? -layer_0[7471-:16] : layer_0[7471-:16]);
                next_layer_0[7487-:16] = (layer_0[7487] ? -layer_0[7487-:16] : layer_0[7487-:16]);
                next_layer_0[7503-:16] = (layer_0[7503] ? -layer_0[7503-:16] : layer_0[7503-:16]);
                next_layer_0[7519-:16] = (layer_0[7519] ? -layer_0[7519-:16] : layer_0[7519-:16]);
                next_layer_0[7535-:16] = (layer_0[7535] ? -layer_0[7535-:16] : layer_0[7535-:16]);
                next_layer_0[7551-:16] = (layer_0[7551] ? -layer_0[7551-:16] : layer_0[7551-:16]);
                next_layer_0[7567-:16] = (layer_0[7567] ? -layer_0[7567-:16] : layer_0[7567-:16]);
                next_layer_0[7583-:16] = (layer_0[7583] ? -layer_0[7583-:16] : layer_0[7583-:16]);
                next_layer_0[7599-:16] = (layer_0[7599] ? -layer_0[7599-:16] : layer_0[7599-:16]);
                next_layer_0[7615-:16] = (layer_0[7615] ? -layer_0[7615-:16] : layer_0[7615-:16]);
                next_layer_0[7631-:16] = (layer_0[7631] ? -layer_0[7631-:16] : layer_0[7631-:16]);
                next_layer_0[7647-:16] = (layer_0[7647] ? -layer_0[7647-:16] : layer_0[7647-:16]);
                next_layer_0[7663-:16] = (layer_0[7663] ? -layer_0[7663-:16] : layer_0[7663-:16]);
                next_layer_0[7679-:16] = (layer_0[7679] ? -layer_0[7679-:16] : layer_0[7679-:16]);
                next_layer_0[7695-:16] = (layer_0[7695] ? -layer_0[7695-:16] : layer_0[7695-:16]);
                next_layer_0[7711-:16] = (layer_0[7711] ? -layer_0[7711-:16] : layer_0[7711-:16]);
                next_layer_0[7727-:16] = (layer_0[7727] ? -layer_0[7727-:16] : layer_0[7727-:16]);
                next_layer_0[7743-:16] = (layer_0[7743] ? -layer_0[7743-:16] : layer_0[7743-:16]);
                next_layer_0[7759-:16] = (layer_0[7759] ? -layer_0[7759-:16] : layer_0[7759-:16]);
                next_layer_0[7775-:16] = (layer_0[7775] ? -layer_0[7775-:16] : layer_0[7775-:16]);
                next_layer_0[7791-:16] = (layer_0[7791] ? -layer_0[7791-:16] : layer_0[7791-:16]);
                next_layer_0[7807-:16] = (layer_0[7807] ? -layer_0[7807-:16] : layer_0[7807-:16]);
                next_layer_0[7823-:16] = (layer_0[7823] ? -layer_0[7823-:16] : layer_0[7823-:16]);
                next_layer_0[7839-:16] = (layer_0[7839] ? -layer_0[7839-:16] : layer_0[7839-:16]);
                next_layer_0[7855-:16] = (layer_0[7855] ? -layer_0[7855-:16] : layer_0[7855-:16]);
                next_layer_0[7871-:16] = (layer_0[7871] ? -layer_0[7871-:16] : layer_0[7871-:16]);
                next_layer_0[7887-:16] = (layer_0[7887] ? -layer_0[7887-:16] : layer_0[7887-:16]);
                next_layer_0[7903-:16] = (layer_0[7903] ? -layer_0[7903-:16] : layer_0[7903-:16]);
                next_layer_0[7919-:16] = (layer_0[7919] ? -layer_0[7919-:16] : layer_0[7919-:16]);
                next_layer_0[7935-:16] = (layer_0[7935] ? -layer_0[7935-:16] : layer_0[7935-:16]);
                next_layer_0[7951-:16] = (layer_0[7951] ? -layer_0[7951-:16] : layer_0[7951-:16]);
                next_layer_0[7967-:16] = (layer_0[7967] ? -layer_0[7967-:16] : layer_0[7967-:16]);
                next_layer_0[7983-:16] = (layer_0[7983] ? -layer_0[7983-:16] : layer_0[7983-:16]);
                next_layer_0[7999-:16] = (layer_0[7999] ? -layer_0[7999-:16] : layer_0[7999-:16]);
                next_layer_0[8015-:16] = (layer_0[8015] ? -layer_0[8015-:16] : layer_0[8015-:16]);
                next_layer_0[8031-:16] = (layer_0[8031] ? -layer_0[8031-:16] : layer_0[8031-:16]);
                next_layer_0[8047-:16] = (layer_0[8047] ? -layer_0[8047-:16] : layer_0[8047-:16]);
                next_layer_0[8063-:16] = (layer_0[8063] ? -layer_0[8063-:16] : layer_0[8063-:16]);
                next_layer_0[8079-:16] = (layer_0[8079] ? -layer_0[8079-:16] : layer_0[8079-:16]);
                next_layer_0[8095-:16] = (layer_0[8095] ? -layer_0[8095-:16] : layer_0[8095-:16]);
                next_layer_0[8111-:16] = (layer_0[8111] ? -layer_0[8111-:16] : layer_0[8111-:16]);
                next_layer_0[8127-:16] = (layer_0[8127] ? -layer_0[8127-:16] : layer_0[8127-:16]);
                next_layer_0[8143-:16] = (layer_0[8143] ? -layer_0[8143-:16] : layer_0[8143-:16]);
                next_layer_0[8159-:16] = (layer_0[8159] ? -layer_0[8159-:16] : layer_0[8159-:16]);
                next_layer_0[8175-:16] = (layer_0[8175] ? -layer_0[8175-:16] : layer_0[8175-:16]);
                next_layer_0[8191-:16] = (layer_0[8191] ? -layer_0[8191-:16] : layer_0[8191-:16]);
                next_layer_0[8207-:16] = (layer_0[8207] ? -layer_0[8207-:16] : layer_0[8207-:16]);
                next_layer_0[8223-:16] = (layer_0[8223] ? -layer_0[8223-:16] : layer_0[8223-:16]);
                next_layer_0[8239-:16] = (layer_0[8239] ? -layer_0[8239-:16] : layer_0[8239-:16]);
                next_layer_0[8255-:16] = (layer_0[8255] ? -layer_0[8255-:16] : layer_0[8255-:16]);
                next_layer_0[8271-:16] = (layer_0[8271] ? -layer_0[8271-:16] : layer_0[8271-:16]);
                next_layer_0[8287-:16] = (layer_0[8287] ? -layer_0[8287-:16] : layer_0[8287-:16]);
                next_layer_0[8303-:16] = (layer_0[8303] ? -layer_0[8303-:16] : layer_0[8303-:16]);
                next_layer_0[8319-:16] = (layer_0[8319] ? -layer_0[8319-:16] : layer_0[8319-:16]);
                next_layer_0[8335-:16] = (layer_0[8335] ? -layer_0[8335-:16] : layer_0[8335-:16]);
                next_layer_0[8351-:16] = (layer_0[8351] ? -layer_0[8351-:16] : layer_0[8351-:16]);
                next_layer_0[8367-:16] = (layer_0[8367] ? -layer_0[8367-:16] : layer_0[8367-:16]);
                next_layer_0[8383-:16] = (layer_0[8383] ? -layer_0[8383-:16] : layer_0[8383-:16]);
                next_layer_0[8399-:16] = (layer_0[8399] ? -layer_0[8399-:16] : layer_0[8399-:16]);
                next_layer_0[8415-:16] = (layer_0[8415] ? -layer_0[8415-:16] : layer_0[8415-:16]);
                next_layer_0[8431-:16] = (layer_0[8431] ? -layer_0[8431-:16] : layer_0[8431-:16]);
                next_layer_0[8447-:16] = (layer_0[8447] ? -layer_0[8447-:16] : layer_0[8447-:16]);
                next_layer_0[8463-:16] = (layer_0[8463] ? -layer_0[8463-:16] : layer_0[8463-:16]);
                next_layer_0[8479-:16] = (layer_0[8479] ? -layer_0[8479-:16] : layer_0[8479-:16]);
                next_layer_0[8495-:16] = (layer_0[8495] ? -layer_0[8495-:16] : layer_0[8495-:16]);
                next_layer_0[8511-:16] = (layer_0[8511] ? -layer_0[8511-:16] : layer_0[8511-:16]);
                next_layer_0[8527-:16] = (layer_0[8527] ? -layer_0[8527-:16] : layer_0[8527-:16]);
                next_layer_0[8543-:16] = (layer_0[8543] ? -layer_0[8543-:16] : layer_0[8543-:16]);
                next_layer_0[8559-:16] = (layer_0[8559] ? -layer_0[8559-:16] : layer_0[8559-:16]);
                next_layer_0[8575-:16] = (layer_0[8575] ? -layer_0[8575-:16] : layer_0[8575-:16]);
                next_layer_0[8591-:16] = (layer_0[8591] ? -layer_0[8591-:16] : layer_0[8591-:16]);
                next_layer_0[8607-:16] = (layer_0[8607] ? -layer_0[8607-:16] : layer_0[8607-:16]);
                next_layer_0[8623-:16] = (layer_0[8623] ? -layer_0[8623-:16] : layer_0[8623-:16]);
                next_layer_0[8639-:16] = (layer_0[8639] ? -layer_0[8639-:16] : layer_0[8639-:16]);
                next_layer_0[8655-:16] = (layer_0[8655] ? -layer_0[8655-:16] : layer_0[8655-:16]);
                next_layer_0[8671-:16] = (layer_0[8671] ? -layer_0[8671-:16] : layer_0[8671-:16]);
                next_layer_0[8687-:16] = (layer_0[8687] ? -layer_0[8687-:16] : layer_0[8687-:16]);
                next_layer_0[8703-:16] = (layer_0[8703] ? -layer_0[8703-:16] : layer_0[8703-:16]);
                next_layer_0[8719-:16] = (layer_0[8719] ? -layer_0[8719-:16] : layer_0[8719-:16]);
                next_layer_0[8735-:16] = (layer_0[8735] ? -layer_0[8735-:16] : layer_0[8735-:16]);
                next_layer_0[8751-:16] = (layer_0[8751] ? -layer_0[8751-:16] : layer_0[8751-:16]);
                next_layer_0[8767-:16] = (layer_0[8767] ? -layer_0[8767-:16] : layer_0[8767-:16]);
                next_layer_0[8783-:16] = (layer_0[8783] ? -layer_0[8783-:16] : layer_0[8783-:16]);
                next_layer_0[8799-:16] = (layer_0[8799] ? -layer_0[8799-:16] : layer_0[8799-:16]);
                next_layer_0[8815-:16] = (layer_0[8815] ? -layer_0[8815-:16] : layer_0[8815-:16]);
                next_layer_0[8831-:16] = (layer_0[8831] ? -layer_0[8831-:16] : layer_0[8831-:16]);
                next_layer_0[8847-:16] = (layer_0[8847] ? -layer_0[8847-:16] : layer_0[8847-:16]);
                next_layer_0[8863-:16] = (layer_0[8863] ? -layer_0[8863-:16] : layer_0[8863-:16]);
                next_layer_0[8879-:16] = (layer_0[8879] ? -layer_0[8879-:16] : layer_0[8879-:16]);
                next_layer_0[8895-:16] = (layer_0[8895] ? -layer_0[8895-:16] : layer_0[8895-:16]);
                next_layer_0[8911-:16] = (layer_0[8911] ? -layer_0[8911-:16] : layer_0[8911-:16]);
                next_layer_0[8927-:16] = (layer_0[8927] ? -layer_0[8927-:16] : layer_0[8927-:16]);
                next_layer_0[8943-:16] = (layer_0[8943] ? -layer_0[8943-:16] : layer_0[8943-:16]);
                next_layer_0[8959-:16] = (layer_0[8959] ? -layer_0[8959-:16] : layer_0[8959-:16]);
                next_layer_0[8975-:16] = (layer_0[8975] ? -layer_0[8975-:16] : layer_0[8975-:16]);
                next_layer_0[8991-:16] = (layer_0[8991] ? -layer_0[8991-:16] : layer_0[8991-:16]);
                next_layer_0[9007-:16] = (layer_0[9007] ? -layer_0[9007-:16] : layer_0[9007-:16]);
                next_layer_0[9023-:16] = (layer_0[9023] ? -layer_0[9023-:16] : layer_0[9023-:16]);
                next_layer_0[9039-:16] = (layer_0[9039] ? -layer_0[9039-:16] : layer_0[9039-:16]);
                next_layer_0[9055-:16] = (layer_0[9055] ? -layer_0[9055-:16] : layer_0[9055-:16]);
                next_layer_0[9071-:16] = (layer_0[9071] ? -layer_0[9071-:16] : layer_0[9071-:16]);
                next_layer_0[9087-:16] = (layer_0[9087] ? -layer_0[9087-:16] : layer_0[9087-:16]);
                next_layer_0[9103-:16] = (layer_0[9103] ? -layer_0[9103-:16] : layer_0[9103-:16]);
                next_layer_0[9119-:16] = (layer_0[9119] ? -layer_0[9119-:16] : layer_0[9119-:16]);
                next_layer_0[9135-:16] = (layer_0[9135] ? -layer_0[9135-:16] : layer_0[9135-:16]);
                next_layer_0[9151-:16] = (layer_0[9151] ? -layer_0[9151-:16] : layer_0[9151-:16]);
                next_layer_0[9167-:16] = (layer_0[9167] ? -layer_0[9167-:16] : layer_0[9167-:16]);
                next_layer_0[9183-:16] = (layer_0[9183] ? -layer_0[9183-:16] : layer_0[9183-:16]);
                next_layer_0[9199-:16] = (layer_0[9199] ? -layer_0[9199-:16] : layer_0[9199-:16]);
                next_layer_0[9215-:16] = (layer_0[9215] ? -layer_0[9215-:16] : layer_0[9215-:16]);
                next_layer_0[9231-:16] = (layer_0[9231] ? -layer_0[9231-:16] : layer_0[9231-:16]);
                next_layer_0[9247-:16] = (layer_0[9247] ? -layer_0[9247-:16] : layer_0[9247-:16]);
                next_layer_0[9263-:16] = (layer_0[9263] ? -layer_0[9263-:16] : layer_0[9263-:16]);
                next_layer_0[9279-:16] = (layer_0[9279] ? -layer_0[9279-:16] : layer_0[9279-:16]);
                next_layer_0[9295-:16] = (layer_0[9295] ? -layer_0[9295-:16] : layer_0[9295-:16]);
                next_layer_0[9311-:16] = (layer_0[9311] ? -layer_0[9311-:16] : layer_0[9311-:16]);
                next_layer_0[9327-:16] = (layer_0[9327] ? -layer_0[9327-:16] : layer_0[9327-:16]);
                next_layer_0[9343-:16] = (layer_0[9343] ? -layer_0[9343-:16] : layer_0[9343-:16]);
                next_layer_0[9359-:16] = (layer_0[9359] ? -layer_0[9359-:16] : layer_0[9359-:16]);
                next_layer_0[9375-:16] = (layer_0[9375] ? -layer_0[9375-:16] : layer_0[9375-:16]);
                next_layer_0[9391-:16] = (layer_0[9391] ? -layer_0[9391-:16] : layer_0[9391-:16]);
                next_layer_0[9407-:16] = (layer_0[9407] ? -layer_0[9407-:16] : layer_0[9407-:16]);
                next_layer_0[9423-:16] = (layer_0[9423] ? -layer_0[9423-:16] : layer_0[9423-:16]);
                next_layer_0[9439-:16] = (layer_0[9439] ? -layer_0[9439-:16] : layer_0[9439-:16]);
                next_layer_0[9455-:16] = (layer_0[9455] ? -layer_0[9455-:16] : layer_0[9455-:16]);
                next_layer_0[9471-:16] = (layer_0[9471] ? -layer_0[9471-:16] : layer_0[9471-:16]);
                next_layer_0[9487-:16] = (layer_0[9487] ? -layer_0[9487-:16] : layer_0[9487-:16]);
                next_layer_0[9503-:16] = (layer_0[9503] ? -layer_0[9503-:16] : layer_0[9503-:16]);
                next_layer_0[9519-:16] = (layer_0[9519] ? -layer_0[9519-:16] : layer_0[9519-:16]);
                next_layer_0[9535-:16] = (layer_0[9535] ? -layer_0[9535-:16] : layer_0[9535-:16]);
                next_layer_0[9551-:16] = (layer_0[9551] ? -layer_0[9551-:16] : layer_0[9551-:16]);
                next_layer_0[9567-:16] = (layer_0[9567] ? -layer_0[9567-:16] : layer_0[9567-:16]);
                next_layer_0[9583-:16] = (layer_0[9583] ? -layer_0[9583-:16] : layer_0[9583-:16]);
                next_layer_0[9599-:16] = (layer_0[9599] ? -layer_0[9599-:16] : layer_0[9599-:16]);
                next_layer_0[9615-:16] = (layer_0[9615] ? -layer_0[9615-:16] : layer_0[9615-:16]);
                next_layer_0[9631-:16] = (layer_0[9631] ? -layer_0[9631-:16] : layer_0[9631-:16]);
                next_layer_0[9647-:16] = (layer_0[9647] ? -layer_0[9647-:16] : layer_0[9647-:16]);
                next_layer_0[9663-:16] = (layer_0[9663] ? -layer_0[9663-:16] : layer_0[9663-:16]);
                next_layer_0[9679-:16] = (layer_0[9679] ? -layer_0[9679-:16] : layer_0[9679-:16]);
                next_layer_0[9695-:16] = (layer_0[9695] ? -layer_0[9695-:16] : layer_0[9695-:16]);
                next_layer_0[9711-:16] = (layer_0[9711] ? -layer_0[9711-:16] : layer_0[9711-:16]);
                next_layer_0[9727-:16] = (layer_0[9727] ? -layer_0[9727-:16] : layer_0[9727-:16]);
                next_layer_0[9743-:16] = (layer_0[9743] ? -layer_0[9743-:16] : layer_0[9743-:16]);
                next_layer_0[9759-:16] = (layer_0[9759] ? -layer_0[9759-:16] : layer_0[9759-:16]);
                next_layer_0[9775-:16] = (layer_0[9775] ? -layer_0[9775-:16] : layer_0[9775-:16]);
                next_layer_0[9791-:16] = (layer_0[9791] ? -layer_0[9791-:16] : layer_0[9791-:16]);
                next_layer_0[9807-:16] = (layer_0[9807] ? -layer_0[9807-:16] : layer_0[9807-:16]);
                next_layer_0[9823-:16] = (layer_0[9823] ? -layer_0[9823-:16] : layer_0[9823-:16]);
                next_layer_0[9839-:16] = (layer_0[9839] ? -layer_0[9839-:16] : layer_0[9839-:16]);
                next_layer_0[9855-:16] = (layer_0[9855] ? -layer_0[9855-:16] : layer_0[9855-:16]);
                next_layer_0[9871-:16] = (layer_0[9871] ? -layer_0[9871-:16] : layer_0[9871-:16]);
                next_layer_0[9887-:16] = (layer_0[9887] ? -layer_0[9887-:16] : layer_0[9887-:16]);
                next_layer_0[9903-:16] = (layer_0[9903] ? -layer_0[9903-:16] : layer_0[9903-:16]);
                next_layer_0[9919-:16] = (layer_0[9919] ? -layer_0[9919-:16] : layer_0[9919-:16]);
                next_layer_0[9935-:16] = (layer_0[9935] ? -layer_0[9935-:16] : layer_0[9935-:16]);
                next_layer_0[9951-:16] = (layer_0[9951] ? -layer_0[9951-:16] : layer_0[9951-:16]);
                next_layer_0[9967-:16] = (layer_0[9967] ? -layer_0[9967-:16] : layer_0[9967-:16]);
                next_layer_0[9983-:16] = (layer_0[9983] ? -layer_0[9983-:16] : layer_0[9983-:16]);
                next_layer_0[9999-:16] = (layer_0[9999] ? -layer_0[9999-:16] : layer_0[9999-:16]);
                next_layer_0[10015-:16] = (layer_0[10015] ? -layer_0[10015-:16] : layer_0[10015-:16]);
                next_layer_0[10031-:16] = (layer_0[10031] ? -layer_0[10031-:16] : layer_0[10031-:16]);
                next_layer_0[10047-:16] = (layer_0[10047] ? -layer_0[10047-:16] : layer_0[10047-:16]);
                next_layer_0[10063-:16] = (layer_0[10063] ? -layer_0[10063-:16] : layer_0[10063-:16]);
                next_layer_0[10079-:16] = (layer_0[10079] ? -layer_0[10079-:16] : layer_0[10079-:16]);
                next_layer_0[10095-:16] = (layer_0[10095] ? -layer_0[10095-:16] : layer_0[10095-:16]);
                next_layer_0[10111-:16] = (layer_0[10111] ? -layer_0[10111-:16] : layer_0[10111-:16]);
                next_layer_0[10127-:16] = (layer_0[10127] ? -layer_0[10127-:16] : layer_0[10127-:16]);
                next_layer_0[10143-:16] = (layer_0[10143] ? -layer_0[10143-:16] : layer_0[10143-:16]);
                next_layer_0[10159-:16] = (layer_0[10159] ? -layer_0[10159-:16] : layer_0[10159-:16]);
                next_layer_0[10175-:16] = (layer_0[10175] ? -layer_0[10175-:16] : layer_0[10175-:16]);
                next_layer_0[10191-:16] = (layer_0[10191] ? -layer_0[10191-:16] : layer_0[10191-:16]);
                next_layer_0[10207-:16] = (layer_0[10207] ? -layer_0[10207-:16] : layer_0[10207-:16]);
                next_layer_0[10223-:16] = (layer_0[10223] ? -layer_0[10223-:16] : layer_0[10223-:16]);
                next_layer_0[10239-:16] = (layer_0[10239] ? -layer_0[10239-:16] : layer_0[10239-:16]);
                next_layer_0[10255-:16] = (layer_0[10255] ? -layer_0[10255-:16] : layer_0[10255-:16]);
                next_layer_0[10271-:16] = (layer_0[10271] ? -layer_0[10271-:16] : layer_0[10271-:16]);
                next_layer_0[10287-:16] = (layer_0[10287] ? -layer_0[10287-:16] : layer_0[10287-:16]);
                next_layer_0[10303-:16] = (layer_0[10303] ? -layer_0[10303-:16] : layer_0[10303-:16]);
                next_layer_0[10319-:16] = (layer_0[10319] ? -layer_0[10319-:16] : layer_0[10319-:16]);
                next_layer_0[10335-:16] = (layer_0[10335] ? -layer_0[10335-:16] : layer_0[10335-:16]);
                next_layer_0[10351-:16] = (layer_0[10351] ? -layer_0[10351-:16] : layer_0[10351-:16]);
                next_layer_0[10367-:16] = (layer_0[10367] ? -layer_0[10367-:16] : layer_0[10367-:16]);
                next_layer_0[10383-:16] = (layer_0[10383] ? -layer_0[10383-:16] : layer_0[10383-:16]);
                next_layer_0[10399-:16] = (layer_0[10399] ? -layer_0[10399-:16] : layer_0[10399-:16]);
                next_layer_0[10415-:16] = (layer_0[10415] ? -layer_0[10415-:16] : layer_0[10415-:16]);
                next_layer_0[10431-:16] = (layer_0[10431] ? -layer_0[10431-:16] : layer_0[10431-:16]);
                next_layer_0[10447-:16] = (layer_0[10447] ? -layer_0[10447-:16] : layer_0[10447-:16]);
                next_layer_0[10463-:16] = (layer_0[10463] ? -layer_0[10463-:16] : layer_0[10463-:16]);
                next_layer_0[10479-:16] = (layer_0[10479] ? -layer_0[10479-:16] : layer_0[10479-:16]);
                next_layer_0[10495-:16] = (layer_0[10495] ? -layer_0[10495-:16] : layer_0[10495-:16]);
                next_layer_0[10511-:16] = (layer_0[10511] ? -layer_0[10511-:16] : layer_0[10511-:16]);
                next_layer_0[10527-:16] = (layer_0[10527] ? -layer_0[10527-:16] : layer_0[10527-:16]);
                next_layer_0[10543-:16] = (layer_0[10543] ? -layer_0[10543-:16] : layer_0[10543-:16]);
                next_layer_0[10559-:16] = (layer_0[10559] ? -layer_0[10559-:16] : layer_0[10559-:16]);
                next_layer_0[10575-:16] = (layer_0[10575] ? -layer_0[10575-:16] : layer_0[10575-:16]);
                next_layer_0[10591-:16] = (layer_0[10591] ? -layer_0[10591-:16] : layer_0[10591-:16]);
                next_layer_0[10607-:16] = (layer_0[10607] ? -layer_0[10607-:16] : layer_0[10607-:16]);
                next_layer_0[10623-:16] = (layer_0[10623] ? -layer_0[10623-:16] : layer_0[10623-:16]);
                next_layer_0[10639-:16] = (layer_0[10639] ? -layer_0[10639-:16] : layer_0[10639-:16]);
                next_layer_0[10655-:16] = (layer_0[10655] ? -layer_0[10655-:16] : layer_0[10655-:16]);
                next_layer_0[10671-:16] = (layer_0[10671] ? -layer_0[10671-:16] : layer_0[10671-:16]);
                next_layer_0[10687-:16] = (layer_0[10687] ? -layer_0[10687-:16] : layer_0[10687-:16]);
                next_layer_0[10703-:16] = (layer_0[10703] ? -layer_0[10703-:16] : layer_0[10703-:16]);
                next_layer_0[10719-:16] = (layer_0[10719] ? -layer_0[10719-:16] : layer_0[10719-:16]);
                next_layer_0[10735-:16] = (layer_0[10735] ? -layer_0[10735-:16] : layer_0[10735-:16]);
                next_layer_0[10751-:16] = (layer_0[10751] ? -layer_0[10751-:16] : layer_0[10751-:16]);
                next_layer_0[10767-:16] = (layer_0[10767] ? -layer_0[10767-:16] : layer_0[10767-:16]);
                next_layer_0[10783-:16] = (layer_0[10783] ? -layer_0[10783-:16] : layer_0[10783-:16]);
                next_layer_0[10799-:16] = (layer_0[10799] ? -layer_0[10799-:16] : layer_0[10799-:16]);
                next_layer_0[10815-:16] = (layer_0[10815] ? -layer_0[10815-:16] : layer_0[10815-:16]);
                next_layer_0[10831-:16] = (layer_0[10831] ? -layer_0[10831-:16] : layer_0[10831-:16]);
                next_layer_0[10847-:16] = (layer_0[10847] ? -layer_0[10847-:16] : layer_0[10847-:16]);
                next_layer_0[10863-:16] = (layer_0[10863] ? -layer_0[10863-:16] : layer_0[10863-:16]);
                next_layer_0[10879-:16] = (layer_0[10879] ? -layer_0[10879-:16] : layer_0[10879-:16]);
                next_layer_0[10895-:16] = (layer_0[10895] ? -layer_0[10895-:16] : layer_0[10895-:16]);
                next_layer_0[10911-:16] = (layer_0[10911] ? -layer_0[10911-:16] : layer_0[10911-:16]);
                next_layer_0[10927-:16] = (layer_0[10927] ? -layer_0[10927-:16] : layer_0[10927-:16]);
                next_layer_0[10943-:16] = (layer_0[10943] ? -layer_0[10943-:16] : layer_0[10943-:16]);
                next_layer_0[10959-:16] = (layer_0[10959] ? -layer_0[10959-:16] : layer_0[10959-:16]);
                next_layer_0[10975-:16] = (layer_0[10975] ? -layer_0[10975-:16] : layer_0[10975-:16]);
                next_layer_0[10991-:16] = (layer_0[10991] ? -layer_0[10991-:16] : layer_0[10991-:16]);
                next_layer_0[11007-:16] = (layer_0[11007] ? -layer_0[11007-:16] : layer_0[11007-:16]);
                next_layer_0[11023-:16] = (layer_0[11023] ? -layer_0[11023-:16] : layer_0[11023-:16]);
                next_layer_0[11039-:16] = (layer_0[11039] ? -layer_0[11039-:16] : layer_0[11039-:16]);
                next_layer_0[11055-:16] = (layer_0[11055] ? -layer_0[11055-:16] : layer_0[11055-:16]);
                next_layer_0[11071-:16] = (layer_0[11071] ? -layer_0[11071-:16] : layer_0[11071-:16]);
                next_layer_0[11087-:16] = (layer_0[11087] ? -layer_0[11087-:16] : layer_0[11087-:16]);
                next_layer_0[11103-:16] = (layer_0[11103] ? -layer_0[11103-:16] : layer_0[11103-:16]);
                next_layer_0[11119-:16] = (layer_0[11119] ? -layer_0[11119-:16] : layer_0[11119-:16]);
                next_layer_0[11135-:16] = (layer_0[11135] ? -layer_0[11135-:16] : layer_0[11135-:16]);
                next_layer_0[11151-:16] = (layer_0[11151] ? -layer_0[11151-:16] : layer_0[11151-:16]);
                next_layer_0[11167-:16] = (layer_0[11167] ? -layer_0[11167-:16] : layer_0[11167-:16]);
                next_layer_0[11183-:16] = (layer_0[11183] ? -layer_0[11183-:16] : layer_0[11183-:16]);
                next_layer_0[11199-:16] = (layer_0[11199] ? -layer_0[11199-:16] : layer_0[11199-:16]);
                next_layer_0[11215-:16] = (layer_0[11215] ? -layer_0[11215-:16] : layer_0[11215-:16]);
                next_layer_0[11231-:16] = (layer_0[11231] ? -layer_0[11231-:16] : layer_0[11231-:16]);
                next_layer_0[11247-:16] = (layer_0[11247] ? -layer_0[11247-:16] : layer_0[11247-:16]);
                next_layer_0[11263-:16] = (layer_0[11263] ? -layer_0[11263-:16] : layer_0[11263-:16]);
                next_layer_0[11279-:16] = (layer_0[11279] ? -layer_0[11279-:16] : layer_0[11279-:16]);
                next_layer_0[11295-:16] = (layer_0[11295] ? -layer_0[11295-:16] : layer_0[11295-:16]);
                next_layer_0[11311-:16] = (layer_0[11311] ? -layer_0[11311-:16] : layer_0[11311-:16]);
                next_layer_0[11327-:16] = (layer_0[11327] ? -layer_0[11327-:16] : layer_0[11327-:16]);
                next_layer_0[11343-:16] = (layer_0[11343] ? -layer_0[11343-:16] : layer_0[11343-:16]);
                next_layer_0[11359-:16] = (layer_0[11359] ? -layer_0[11359-:16] : layer_0[11359-:16]);
                next_layer_0[11375-:16] = (layer_0[11375] ? -layer_0[11375-:16] : layer_0[11375-:16]);
                next_layer_0[11391-:16] = (layer_0[11391] ? -layer_0[11391-:16] : layer_0[11391-:16]);
                next_layer_0[11407-:16] = (layer_0[11407] ? -layer_0[11407-:16] : layer_0[11407-:16]);
                next_layer_0[11423-:16] = (layer_0[11423] ? -layer_0[11423-:16] : layer_0[11423-:16]);
                next_layer_0[11439-:16] = (layer_0[11439] ? -layer_0[11439-:16] : layer_0[11439-:16]);
                next_layer_0[11455-:16] = (layer_0[11455] ? -layer_0[11455-:16] : layer_0[11455-:16]);
                next_layer_0[11471-:16] = (layer_0[11471] ? -layer_0[11471-:16] : layer_0[11471-:16]);
                next_layer_0[11487-:16] = (layer_0[11487] ? -layer_0[11487-:16] : layer_0[11487-:16]);
                next_layer_0[11503-:16] = (layer_0[11503] ? -layer_0[11503-:16] : layer_0[11503-:16]);
                next_layer_0[11519-:16] = (layer_0[11519] ? -layer_0[11519-:16] : layer_0[11519-:16]);
                next_layer_0[11535-:16] = (layer_0[11535] ? -layer_0[11535-:16] : layer_0[11535-:16]);
                next_layer_0[11551-:16] = (layer_0[11551] ? -layer_0[11551-:16] : layer_0[11551-:16]);
                next_layer_0[11567-:16] = (layer_0[11567] ? -layer_0[11567-:16] : layer_0[11567-:16]);
                next_layer_0[11583-:16] = (layer_0[11583] ? -layer_0[11583-:16] : layer_0[11583-:16]);
                next_layer_0[11599-:16] = (layer_0[11599] ? -layer_0[11599-:16] : layer_0[11599-:16]);
                next_layer_0[11615-:16] = (layer_0[11615] ? -layer_0[11615-:16] : layer_0[11615-:16]);
                next_layer_0[11631-:16] = (layer_0[11631] ? -layer_0[11631-:16] : layer_0[11631-:16]);
                next_layer_0[11647-:16] = (layer_0[11647] ? -layer_0[11647-:16] : layer_0[11647-:16]);
                next_layer_0[11663-:16] = (layer_0[11663] ? -layer_0[11663-:16] : layer_0[11663-:16]);
                next_layer_0[11679-:16] = (layer_0[11679] ? -layer_0[11679-:16] : layer_0[11679-:16]);
                next_layer_0[11695-:16] = (layer_0[11695] ? -layer_0[11695-:16] : layer_0[11695-:16]);
                next_layer_0[11711-:16] = (layer_0[11711] ? -layer_0[11711-:16] : layer_0[11711-:16]);
                next_layer_0[11727-:16] = (layer_0[11727] ? -layer_0[11727-:16] : layer_0[11727-:16]);
                next_layer_0[11743-:16] = (layer_0[11743] ? -layer_0[11743-:16] : layer_0[11743-:16]);
                next_layer_0[11759-:16] = (layer_0[11759] ? -layer_0[11759-:16] : layer_0[11759-:16]);
                next_layer_0[11775-:16] = (layer_0[11775] ? -layer_0[11775-:16] : layer_0[11775-:16]);
                next_layer_0[11791-:16] = (layer_0[11791] ? -layer_0[11791-:16] : layer_0[11791-:16]);
                next_layer_0[11807-:16] = (layer_0[11807] ? -layer_0[11807-:16] : layer_0[11807-:16]);
                next_layer_0[11823-:16] = (layer_0[11823] ? -layer_0[11823-:16] : layer_0[11823-:16]);
                next_layer_0[11839-:16] = (layer_0[11839] ? -layer_0[11839-:16] : layer_0[11839-:16]);
                next_layer_0[11855-:16] = (layer_0[11855] ? -layer_0[11855-:16] : layer_0[11855-:16]);
                next_layer_0[11871-:16] = (layer_0[11871] ? -layer_0[11871-:16] : layer_0[11871-:16]);
                next_layer_0[11887-:16] = (layer_0[11887] ? -layer_0[11887-:16] : layer_0[11887-:16]);
                next_layer_0[11903-:16] = (layer_0[11903] ? -layer_0[11903-:16] : layer_0[11903-:16]);
                next_layer_0[11919-:16] = (layer_0[11919] ? -layer_0[11919-:16] : layer_0[11919-:16]);
                next_layer_0[11935-:16] = (layer_0[11935] ? -layer_0[11935-:16] : layer_0[11935-:16]);
                next_layer_0[11951-:16] = (layer_0[11951] ? -layer_0[11951-:16] : layer_0[11951-:16]);
                next_layer_0[11967-:16] = (layer_0[11967] ? -layer_0[11967-:16] : layer_0[11967-:16]);
                next_layer_0[11983-:16] = (layer_0[11983] ? -layer_0[11983-:16] : layer_0[11983-:16]);
                next_layer_0[11999-:16] = (layer_0[11999] ? -layer_0[11999-:16] : layer_0[11999-:16]);
                next_layer_0[12015-:16] = (layer_0[12015] ? -layer_0[12015-:16] : layer_0[12015-:16]);
                next_layer_0[12031-:16] = (layer_0[12031] ? -layer_0[12031-:16] : layer_0[12031-:16]);
                next_layer_0[12047-:16] = (layer_0[12047] ? -layer_0[12047-:16] : layer_0[12047-:16]);
                next_layer_0[12063-:16] = (layer_0[12063] ? -layer_0[12063-:16] : layer_0[12063-:16]);
                next_layer_0[12079-:16] = (layer_0[12079] ? -layer_0[12079-:16] : layer_0[12079-:16]);
                next_layer_0[12095-:16] = (layer_0[12095] ? -layer_0[12095-:16] : layer_0[12095-:16]);
                next_layer_0[12111-:16] = (layer_0[12111] ? -layer_0[12111-:16] : layer_0[12111-:16]);
                next_layer_0[12127-:16] = (layer_0[12127] ? -layer_0[12127-:16] : layer_0[12127-:16]);
                next_layer_0[12143-:16] = (layer_0[12143] ? -layer_0[12143-:16] : layer_0[12143-:16]);
                next_layer_0[12159-:16] = (layer_0[12159] ? -layer_0[12159-:16] : layer_0[12159-:16]);
                next_layer_0[12175-:16] = (layer_0[12175] ? -layer_0[12175-:16] : layer_0[12175-:16]);
                next_layer_0[12191-:16] = (layer_0[12191] ? -layer_0[12191-:16] : layer_0[12191-:16]);
                next_layer_0[12207-:16] = (layer_0[12207] ? -layer_0[12207-:16] : layer_0[12207-:16]);
                next_layer_0[12223-:16] = (layer_0[12223] ? -layer_0[12223-:16] : layer_0[12223-:16]);
                next_layer_0[12239-:16] = (layer_0[12239] ? -layer_0[12239-:16] : layer_0[12239-:16]);
                next_layer_0[12255-:16] = (layer_0[12255] ? -layer_0[12255-:16] : layer_0[12255-:16]);
                next_layer_0[12271-:16] = (layer_0[12271] ? -layer_0[12271-:16] : layer_0[12271-:16]);
                next_layer_0[12287-:16] = (layer_0[12287] ? -layer_0[12287-:16] : layer_0[12287-:16]);
                next_layer_0[12303-:16] = (layer_0[12303] ? -layer_0[12303-:16] : layer_0[12303-:16]);
                next_layer_0[12319-:16] = (layer_0[12319] ? -layer_0[12319-:16] : layer_0[12319-:16]);
                next_layer_0[12335-:16] = (layer_0[12335] ? -layer_0[12335-:16] : layer_0[12335-:16]);
                next_layer_0[12351-:16] = (layer_0[12351] ? -layer_0[12351-:16] : layer_0[12351-:16]);
                next_layer_0[12367-:16] = (layer_0[12367] ? -layer_0[12367-:16] : layer_0[12367-:16]);
                next_layer_0[12383-:16] = (layer_0[12383] ? -layer_0[12383-:16] : layer_0[12383-:16]);
                next_layer_0[12399-:16] = (layer_0[12399] ? -layer_0[12399-:16] : layer_0[12399-:16]);
                next_layer_0[12415-:16] = (layer_0[12415] ? -layer_0[12415-:16] : layer_0[12415-:16]);
                next_layer_0[12431-:16] = (layer_0[12431] ? -layer_0[12431-:16] : layer_0[12431-:16]);
                next_layer_0[12447-:16] = (layer_0[12447] ? -layer_0[12447-:16] : layer_0[12447-:16]);
                next_layer_0[12463-:16] = (layer_0[12463] ? -layer_0[12463-:16] : layer_0[12463-:16]);
                next_layer_0[12479-:16] = (layer_0[12479] ? -layer_0[12479-:16] : layer_0[12479-:16]);
                next_layer_0[12495-:16] = (layer_0[12495] ? -layer_0[12495-:16] : layer_0[12495-:16]);
                next_layer_0[12511-:16] = (layer_0[12511] ? -layer_0[12511-:16] : layer_0[12511-:16]);
                next_layer_0[12527-:16] = (layer_0[12527] ? -layer_0[12527-:16] : layer_0[12527-:16]);
                next_layer_0[12543-:16] = (layer_0[12543] ? -layer_0[12543-:16] : layer_0[12543-:16]);
            end
            SBIAS: begin
                next_layer_0[15-:16] = layer_0[15-:16] + bias_0[15-:16];
                next_layer_0[31-:16] = layer_0[31-:16] + bias_0[31-:16];
                next_layer_0[47-:16] = layer_0[47-:16] + bias_0[47-:16];
                next_layer_0[63-:16] = layer_0[63-:16] + bias_0[63-:16];
                next_layer_0[79-:16] = layer_0[79-:16] + bias_0[79-:16];
                next_layer_0[95-:16] = layer_0[95-:16] + bias_0[95-:16];
                next_layer_0[111-:16] = layer_0[111-:16] + bias_0[111-:16];
                next_layer_0[127-:16] = layer_0[127-:16] + bias_0[127-:16];
                next_layer_0[143-:16] = layer_0[143-:16] + bias_0[143-:16];
                next_layer_0[159-:16] = layer_0[159-:16] + bias_0[159-:16];
                next_layer_0[175-:16] = layer_0[175-:16] + bias_0[175-:16];
                next_layer_0[191-:16] = layer_0[191-:16] + bias_0[191-:16];
                next_layer_0[207-:16] = layer_0[207-:16] + bias_0[207-:16];
                next_layer_0[223-:16] = layer_0[223-:16] + bias_0[223-:16];
                next_layer_0[239-:16] = layer_0[239-:16] + bias_0[239-:16];
                next_layer_0[255-:16] = layer_0[255-:16] + bias_0[255-:16];
                next_layer_0[271-:16] = layer_0[271-:16] + bias_0[271-:16];
                next_layer_0[287-:16] = layer_0[287-:16] + bias_0[287-:16];
                next_layer_0[303-:16] = layer_0[303-:16] + bias_0[303-:16];
                next_layer_0[319-:16] = layer_0[319-:16] + bias_0[319-:16];
                next_layer_0[335-:16] = layer_0[335-:16] + bias_0[335-:16];
                next_layer_0[351-:16] = layer_0[351-:16] + bias_0[351-:16];
                next_layer_0[367-:16] = layer_0[367-:16] + bias_0[367-:16];
                next_layer_0[383-:16] = layer_0[383-:16] + bias_0[383-:16];
                next_layer_0[399-:16] = layer_0[399-:16] + bias_0[399-:16];
                next_layer_0[415-:16] = layer_0[415-:16] + bias_0[415-:16];
                next_layer_0[431-:16] = layer_0[431-:16] + bias_0[431-:16];
                next_layer_0[447-:16] = layer_0[447-:16] + bias_0[447-:16];
                next_layer_0[463-:16] = layer_0[463-:16] + bias_0[463-:16];
                next_layer_0[479-:16] = layer_0[479-:16] + bias_0[479-:16];
                next_layer_0[495-:16] = layer_0[495-:16] + bias_0[495-:16];
                next_layer_0[511-:16] = layer_0[511-:16] + bias_0[511-:16];
                next_layer_0[527-:16] = layer_0[527-:16] + bias_0[527-:16];
                next_layer_0[543-:16] = layer_0[543-:16] + bias_0[543-:16];
                next_layer_0[559-:16] = layer_0[559-:16] + bias_0[559-:16];
                next_layer_0[575-:16] = layer_0[575-:16] + bias_0[575-:16];
                next_layer_0[591-:16] = layer_0[591-:16] + bias_0[591-:16];
                next_layer_0[607-:16] = layer_0[607-:16] + bias_0[607-:16];
                next_layer_0[623-:16] = layer_0[623-:16] + bias_0[623-:16];
                next_layer_0[639-:16] = layer_0[639-:16] + bias_0[639-:16];
                next_layer_0[655-:16] = layer_0[655-:16] + bias_0[655-:16];
                next_layer_0[671-:16] = layer_0[671-:16] + bias_0[671-:16];
                next_layer_0[687-:16] = layer_0[687-:16] + bias_0[687-:16];
                next_layer_0[703-:16] = layer_0[703-:16] + bias_0[703-:16];
                next_layer_0[719-:16] = layer_0[719-:16] + bias_0[719-:16];
                next_layer_0[735-:16] = layer_0[735-:16] + bias_0[735-:16];
                next_layer_0[751-:16] = layer_0[751-:16] + bias_0[751-:16];
                next_layer_0[767-:16] = layer_0[767-:16] + bias_0[767-:16];
                next_layer_0[783-:16] = layer_0[783-:16] + bias_0[783-:16];
                next_layer_0[799-:16] = layer_0[799-:16] + bias_0[799-:16];
                next_layer_0[815-:16] = layer_0[815-:16] + bias_0[815-:16];
                next_layer_0[831-:16] = layer_0[831-:16] + bias_0[831-:16];
                next_layer_0[847-:16] = layer_0[847-:16] + bias_0[847-:16];
                next_layer_0[863-:16] = layer_0[863-:16] + bias_0[863-:16];
                next_layer_0[879-:16] = layer_0[879-:16] + bias_0[879-:16];
                next_layer_0[895-:16] = layer_0[895-:16] + bias_0[895-:16];
                next_layer_0[911-:16] = layer_0[911-:16] + bias_0[911-:16];
                next_layer_0[927-:16] = layer_0[927-:16] + bias_0[927-:16];
                next_layer_0[943-:16] = layer_0[943-:16] + bias_0[943-:16];
                next_layer_0[959-:16] = layer_0[959-:16] + bias_0[959-:16];
                next_layer_0[975-:16] = layer_0[975-:16] + bias_0[975-:16];
                next_layer_0[991-:16] = layer_0[991-:16] + bias_0[991-:16];
                next_layer_0[1007-:16] = layer_0[1007-:16] + bias_0[1007-:16];
                next_layer_0[1023-:16] = layer_0[1023-:16] + bias_0[1023-:16];
                next_layer_0[1039-:16] = layer_0[1039-:16] + bias_0[1039-:16];
                next_layer_0[1055-:16] = layer_0[1055-:16] + bias_0[1055-:16];
                next_layer_0[1071-:16] = layer_0[1071-:16] + bias_0[1071-:16];
                next_layer_0[1087-:16] = layer_0[1087-:16] + bias_0[1087-:16];
                next_layer_0[1103-:16] = layer_0[1103-:16] + bias_0[1103-:16];
                next_layer_0[1119-:16] = layer_0[1119-:16] + bias_0[1119-:16];
                next_layer_0[1135-:16] = layer_0[1135-:16] + bias_0[1135-:16];
                next_layer_0[1151-:16] = layer_0[1151-:16] + bias_0[1151-:16];
                next_layer_0[1167-:16] = layer_0[1167-:16] + bias_0[1167-:16];
                next_layer_0[1183-:16] = layer_0[1183-:16] + bias_0[1183-:16];
                next_layer_0[1199-:16] = layer_0[1199-:16] + bias_0[1199-:16];
                next_layer_0[1215-:16] = layer_0[1215-:16] + bias_0[1215-:16];
                next_layer_0[1231-:16] = layer_0[1231-:16] + bias_0[1231-:16];
                next_layer_0[1247-:16] = layer_0[1247-:16] + bias_0[1247-:16];
                next_layer_0[1263-:16] = layer_0[1263-:16] + bias_0[1263-:16];
                next_layer_0[1279-:16] = layer_0[1279-:16] + bias_0[1279-:16];
                next_layer_0[1295-:16] = layer_0[1295-:16] + bias_0[1295-:16];
                next_layer_0[1311-:16] = layer_0[1311-:16] + bias_0[1311-:16];
                next_layer_0[1327-:16] = layer_0[1327-:16] + bias_0[1327-:16];
                next_layer_0[1343-:16] = layer_0[1343-:16] + bias_0[1343-:16];
                next_layer_0[1359-:16] = layer_0[1359-:16] + bias_0[1359-:16];
                next_layer_0[1375-:16] = layer_0[1375-:16] + bias_0[1375-:16];
                next_layer_0[1391-:16] = layer_0[1391-:16] + bias_0[1391-:16];
                next_layer_0[1407-:16] = layer_0[1407-:16] + bias_0[1407-:16];
                next_layer_0[1423-:16] = layer_0[1423-:16] + bias_0[1423-:16];
                next_layer_0[1439-:16] = layer_0[1439-:16] + bias_0[1439-:16];
                next_layer_0[1455-:16] = layer_0[1455-:16] + bias_0[1455-:16];
                next_layer_0[1471-:16] = layer_0[1471-:16] + bias_0[1471-:16];
                next_layer_0[1487-:16] = layer_0[1487-:16] + bias_0[1487-:16];
                next_layer_0[1503-:16] = layer_0[1503-:16] + bias_0[1503-:16];
                next_layer_0[1519-:16] = layer_0[1519-:16] + bias_0[1519-:16];
                next_layer_0[1535-:16] = layer_0[1535-:16] + bias_0[1535-:16];
                next_layer_0[1551-:16] = layer_0[1551-:16] + bias_0[1551-:16];
                next_layer_0[1567-:16] = layer_0[1567-:16] + bias_0[1567-:16];
                next_layer_0[1583-:16] = layer_0[1583-:16] + bias_0[1583-:16];
                next_layer_0[1599-:16] = layer_0[1599-:16] + bias_0[1599-:16];
                next_layer_0[1615-:16] = layer_0[1615-:16] + bias_0[1615-:16];
                next_layer_0[1631-:16] = layer_0[1631-:16] + bias_0[1631-:16];
                next_layer_0[1647-:16] = layer_0[1647-:16] + bias_0[1647-:16];
                next_layer_0[1663-:16] = layer_0[1663-:16] + bias_0[1663-:16];
                next_layer_0[1679-:16] = layer_0[1679-:16] + bias_0[1679-:16];
                next_layer_0[1695-:16] = layer_0[1695-:16] + bias_0[1695-:16];
                next_layer_0[1711-:16] = layer_0[1711-:16] + bias_0[1711-:16];
                next_layer_0[1727-:16] = layer_0[1727-:16] + bias_0[1727-:16];
                next_layer_0[1743-:16] = layer_0[1743-:16] + bias_0[1743-:16];
                next_layer_0[1759-:16] = layer_0[1759-:16] + bias_0[1759-:16];
                next_layer_0[1775-:16] = layer_0[1775-:16] + bias_0[1775-:16];
                next_layer_0[1791-:16] = layer_0[1791-:16] + bias_0[1791-:16];
                next_layer_0[1807-:16] = layer_0[1807-:16] + bias_0[1807-:16];
                next_layer_0[1823-:16] = layer_0[1823-:16] + bias_0[1823-:16];
                next_layer_0[1839-:16] = layer_0[1839-:16] + bias_0[1839-:16];
                next_layer_0[1855-:16] = layer_0[1855-:16] + bias_0[1855-:16];
                next_layer_0[1871-:16] = layer_0[1871-:16] + bias_0[1871-:16];
                next_layer_0[1887-:16] = layer_0[1887-:16] + bias_0[1887-:16];
                next_layer_0[1903-:16] = layer_0[1903-:16] + bias_0[1903-:16];
                next_layer_0[1919-:16] = layer_0[1919-:16] + bias_0[1919-:16];
                next_layer_0[1935-:16] = layer_0[1935-:16] + bias_0[1935-:16];
                next_layer_0[1951-:16] = layer_0[1951-:16] + bias_0[1951-:16];
                next_layer_0[1967-:16] = layer_0[1967-:16] + bias_0[1967-:16];
                next_layer_0[1983-:16] = layer_0[1983-:16] + bias_0[1983-:16];
                next_layer_0[1999-:16] = layer_0[1999-:16] + bias_0[1999-:16];
                next_layer_0[2015-:16] = layer_0[2015-:16] + bias_0[2015-:16];
                next_layer_0[2031-:16] = layer_0[2031-:16] + bias_0[2031-:16];
                next_layer_0[2047-:16] = layer_0[2047-:16] + bias_0[2047-:16];
                next_layer_0[2063-:16] = layer_0[2063-:16] + bias_0[2063-:16];
                next_layer_0[2079-:16] = layer_0[2079-:16] + bias_0[2079-:16];
                next_layer_0[2095-:16] = layer_0[2095-:16] + bias_0[2095-:16];
                next_layer_0[2111-:16] = layer_0[2111-:16] + bias_0[2111-:16];
                next_layer_0[2127-:16] = layer_0[2127-:16] + bias_0[2127-:16];
                next_layer_0[2143-:16] = layer_0[2143-:16] + bias_0[2143-:16];
                next_layer_0[2159-:16] = layer_0[2159-:16] + bias_0[2159-:16];
                next_layer_0[2175-:16] = layer_0[2175-:16] + bias_0[2175-:16];
                next_layer_0[2191-:16] = layer_0[2191-:16] + bias_0[2191-:16];
                next_layer_0[2207-:16] = layer_0[2207-:16] + bias_0[2207-:16];
                next_layer_0[2223-:16] = layer_0[2223-:16] + bias_0[2223-:16];
                next_layer_0[2239-:16] = layer_0[2239-:16] + bias_0[2239-:16];
                next_layer_0[2255-:16] = layer_0[2255-:16] + bias_0[2255-:16];
                next_layer_0[2271-:16] = layer_0[2271-:16] + bias_0[2271-:16];
                next_layer_0[2287-:16] = layer_0[2287-:16] + bias_0[2287-:16];
                next_layer_0[2303-:16] = layer_0[2303-:16] + bias_0[2303-:16];
                next_layer_0[2319-:16] = layer_0[2319-:16] + bias_0[2319-:16];
                next_layer_0[2335-:16] = layer_0[2335-:16] + bias_0[2335-:16];
                next_layer_0[2351-:16] = layer_0[2351-:16] + bias_0[2351-:16];
                next_layer_0[2367-:16] = layer_0[2367-:16] + bias_0[2367-:16];
                next_layer_0[2383-:16] = layer_0[2383-:16] + bias_0[2383-:16];
                next_layer_0[2399-:16] = layer_0[2399-:16] + bias_0[2399-:16];
                next_layer_0[2415-:16] = layer_0[2415-:16] + bias_0[2415-:16];
                next_layer_0[2431-:16] = layer_0[2431-:16] + bias_0[2431-:16];
                next_layer_0[2447-:16] = layer_0[2447-:16] + bias_0[2447-:16];
                next_layer_0[2463-:16] = layer_0[2463-:16] + bias_0[2463-:16];
                next_layer_0[2479-:16] = layer_0[2479-:16] + bias_0[2479-:16];
                next_layer_0[2495-:16] = layer_0[2495-:16] + bias_0[2495-:16];
                next_layer_0[2511-:16] = layer_0[2511-:16] + bias_0[2511-:16];
                next_layer_0[2527-:16] = layer_0[2527-:16] + bias_0[2527-:16];
                next_layer_0[2543-:16] = layer_0[2543-:16] + bias_0[2543-:16];
                next_layer_0[2559-:16] = layer_0[2559-:16] + bias_0[2559-:16];
                next_layer_0[2575-:16] = layer_0[2575-:16] + bias_0[2575-:16];
                next_layer_0[2591-:16] = layer_0[2591-:16] + bias_0[2591-:16];
                next_layer_0[2607-:16] = layer_0[2607-:16] + bias_0[2607-:16];
                next_layer_0[2623-:16] = layer_0[2623-:16] + bias_0[2623-:16];
                next_layer_0[2639-:16] = layer_0[2639-:16] + bias_0[2639-:16];
                next_layer_0[2655-:16] = layer_0[2655-:16] + bias_0[2655-:16];
                next_layer_0[2671-:16] = layer_0[2671-:16] + bias_0[2671-:16];
                next_layer_0[2687-:16] = layer_0[2687-:16] + bias_0[2687-:16];
                next_layer_0[2703-:16] = layer_0[2703-:16] + bias_0[2703-:16];
                next_layer_0[2719-:16] = layer_0[2719-:16] + bias_0[2719-:16];
                next_layer_0[2735-:16] = layer_0[2735-:16] + bias_0[2735-:16];
                next_layer_0[2751-:16] = layer_0[2751-:16] + bias_0[2751-:16];
                next_layer_0[2767-:16] = layer_0[2767-:16] + bias_0[2767-:16];
                next_layer_0[2783-:16] = layer_0[2783-:16] + bias_0[2783-:16];
                next_layer_0[2799-:16] = layer_0[2799-:16] + bias_0[2799-:16];
                next_layer_0[2815-:16] = layer_0[2815-:16] + bias_0[2815-:16];
                next_layer_0[2831-:16] = layer_0[2831-:16] + bias_0[2831-:16];
                next_layer_0[2847-:16] = layer_0[2847-:16] + bias_0[2847-:16];
                next_layer_0[2863-:16] = layer_0[2863-:16] + bias_0[2863-:16];
                next_layer_0[2879-:16] = layer_0[2879-:16] + bias_0[2879-:16];
                next_layer_0[2895-:16] = layer_0[2895-:16] + bias_0[2895-:16];
                next_layer_0[2911-:16] = layer_0[2911-:16] + bias_0[2911-:16];
                next_layer_0[2927-:16] = layer_0[2927-:16] + bias_0[2927-:16];
                next_layer_0[2943-:16] = layer_0[2943-:16] + bias_0[2943-:16];
                next_layer_0[2959-:16] = layer_0[2959-:16] + bias_0[2959-:16];
                next_layer_0[2975-:16] = layer_0[2975-:16] + bias_0[2975-:16];
                next_layer_0[2991-:16] = layer_0[2991-:16] + bias_0[2991-:16];
                next_layer_0[3007-:16] = layer_0[3007-:16] + bias_0[3007-:16];
                next_layer_0[3023-:16] = layer_0[3023-:16] + bias_0[3023-:16];
                next_layer_0[3039-:16] = layer_0[3039-:16] + bias_0[3039-:16];
                next_layer_0[3055-:16] = layer_0[3055-:16] + bias_0[3055-:16];
                next_layer_0[3071-:16] = layer_0[3071-:16] + bias_0[3071-:16];
                next_layer_0[3087-:16] = layer_0[3087-:16] + bias_0[3087-:16];
                next_layer_0[3103-:16] = layer_0[3103-:16] + bias_0[3103-:16];
                next_layer_0[3119-:16] = layer_0[3119-:16] + bias_0[3119-:16];
                next_layer_0[3135-:16] = layer_0[3135-:16] + bias_0[3135-:16];
                next_layer_0[3151-:16] = layer_0[3151-:16] + bias_0[3151-:16];
                next_layer_0[3167-:16] = layer_0[3167-:16] + bias_0[3167-:16];
                next_layer_0[3183-:16] = layer_0[3183-:16] + bias_0[3183-:16];
                next_layer_0[3199-:16] = layer_0[3199-:16] + bias_0[3199-:16];
                next_layer_0[3215-:16] = layer_0[3215-:16] + bias_0[3215-:16];
                next_layer_0[3231-:16] = layer_0[3231-:16] + bias_0[3231-:16];
                next_layer_0[3247-:16] = layer_0[3247-:16] + bias_0[3247-:16];
                next_layer_0[3263-:16] = layer_0[3263-:16] + bias_0[3263-:16];
                next_layer_0[3279-:16] = layer_0[3279-:16] + bias_0[3279-:16];
                next_layer_0[3295-:16] = layer_0[3295-:16] + bias_0[3295-:16];
                next_layer_0[3311-:16] = layer_0[3311-:16] + bias_0[3311-:16];
                next_layer_0[3327-:16] = layer_0[3327-:16] + bias_0[3327-:16];
                next_layer_0[3343-:16] = layer_0[3343-:16] + bias_0[3343-:16];
                next_layer_0[3359-:16] = layer_0[3359-:16] + bias_0[3359-:16];
                next_layer_0[3375-:16] = layer_0[3375-:16] + bias_0[3375-:16];
                next_layer_0[3391-:16] = layer_0[3391-:16] + bias_0[3391-:16];
                next_layer_0[3407-:16] = layer_0[3407-:16] + bias_0[3407-:16];
                next_layer_0[3423-:16] = layer_0[3423-:16] + bias_0[3423-:16];
                next_layer_0[3439-:16] = layer_0[3439-:16] + bias_0[3439-:16];
                next_layer_0[3455-:16] = layer_0[3455-:16] + bias_0[3455-:16];
                next_layer_0[3471-:16] = layer_0[3471-:16] + bias_0[3471-:16];
                next_layer_0[3487-:16] = layer_0[3487-:16] + bias_0[3487-:16];
                next_layer_0[3503-:16] = layer_0[3503-:16] + bias_0[3503-:16];
                next_layer_0[3519-:16] = layer_0[3519-:16] + bias_0[3519-:16];
                next_layer_0[3535-:16] = layer_0[3535-:16] + bias_0[3535-:16];
                next_layer_0[3551-:16] = layer_0[3551-:16] + bias_0[3551-:16];
                next_layer_0[3567-:16] = layer_0[3567-:16] + bias_0[3567-:16];
                next_layer_0[3583-:16] = layer_0[3583-:16] + bias_0[3583-:16];
                next_layer_0[3599-:16] = layer_0[3599-:16] + bias_0[3599-:16];
                next_layer_0[3615-:16] = layer_0[3615-:16] + bias_0[3615-:16];
                next_layer_0[3631-:16] = layer_0[3631-:16] + bias_0[3631-:16];
                next_layer_0[3647-:16] = layer_0[3647-:16] + bias_0[3647-:16];
                next_layer_0[3663-:16] = layer_0[3663-:16] + bias_0[3663-:16];
                next_layer_0[3679-:16] = layer_0[3679-:16] + bias_0[3679-:16];
                next_layer_0[3695-:16] = layer_0[3695-:16] + bias_0[3695-:16];
                next_layer_0[3711-:16] = layer_0[3711-:16] + bias_0[3711-:16];
                next_layer_0[3727-:16] = layer_0[3727-:16] + bias_0[3727-:16];
                next_layer_0[3743-:16] = layer_0[3743-:16] + bias_0[3743-:16];
                next_layer_0[3759-:16] = layer_0[3759-:16] + bias_0[3759-:16];
                next_layer_0[3775-:16] = layer_0[3775-:16] + bias_0[3775-:16];
                next_layer_0[3791-:16] = layer_0[3791-:16] + bias_0[3791-:16];
                next_layer_0[3807-:16] = layer_0[3807-:16] + bias_0[3807-:16];
                next_layer_0[3823-:16] = layer_0[3823-:16] + bias_0[3823-:16];
                next_layer_0[3839-:16] = layer_0[3839-:16] + bias_0[3839-:16];
                next_layer_0[3855-:16] = layer_0[3855-:16] + bias_0[3855-:16];
                next_layer_0[3871-:16] = layer_0[3871-:16] + bias_0[3871-:16];
                next_layer_0[3887-:16] = layer_0[3887-:16] + bias_0[3887-:16];
                next_layer_0[3903-:16] = layer_0[3903-:16] + bias_0[3903-:16];
                next_layer_0[3919-:16] = layer_0[3919-:16] + bias_0[3919-:16];
                next_layer_0[3935-:16] = layer_0[3935-:16] + bias_0[3935-:16];
                next_layer_0[3951-:16] = layer_0[3951-:16] + bias_0[3951-:16];
                next_layer_0[3967-:16] = layer_0[3967-:16] + bias_0[3967-:16];
                next_layer_0[3983-:16] = layer_0[3983-:16] + bias_0[3983-:16];
                next_layer_0[3999-:16] = layer_0[3999-:16] + bias_0[3999-:16];
                next_layer_0[4015-:16] = layer_0[4015-:16] + bias_0[4015-:16];
                next_layer_0[4031-:16] = layer_0[4031-:16] + bias_0[4031-:16];
                next_layer_0[4047-:16] = layer_0[4047-:16] + bias_0[4047-:16];
                next_layer_0[4063-:16] = layer_0[4063-:16] + bias_0[4063-:16];
                next_layer_0[4079-:16] = layer_0[4079-:16] + bias_0[4079-:16];
                next_layer_0[4095-:16] = layer_0[4095-:16] + bias_0[4095-:16];
                next_layer_0[4111-:16] = layer_0[4111-:16] + bias_0[4111-:16];
                next_layer_0[4127-:16] = layer_0[4127-:16] + bias_0[4127-:16];
                next_layer_0[4143-:16] = layer_0[4143-:16] + bias_0[4143-:16];
                next_layer_0[4159-:16] = layer_0[4159-:16] + bias_0[4159-:16];
                next_layer_0[4175-:16] = layer_0[4175-:16] + bias_0[4175-:16];
                next_layer_0[4191-:16] = layer_0[4191-:16] + bias_0[4191-:16];
                next_layer_0[4207-:16] = layer_0[4207-:16] + bias_0[4207-:16];
                next_layer_0[4223-:16] = layer_0[4223-:16] + bias_0[4223-:16];
                next_layer_0[4239-:16] = layer_0[4239-:16] + bias_0[4239-:16];
                next_layer_0[4255-:16] = layer_0[4255-:16] + bias_0[4255-:16];
                next_layer_0[4271-:16] = layer_0[4271-:16] + bias_0[4271-:16];
                next_layer_0[4287-:16] = layer_0[4287-:16] + bias_0[4287-:16];
                next_layer_0[4303-:16] = layer_0[4303-:16] + bias_0[4303-:16];
                next_layer_0[4319-:16] = layer_0[4319-:16] + bias_0[4319-:16];
                next_layer_0[4335-:16] = layer_0[4335-:16] + bias_0[4335-:16];
                next_layer_0[4351-:16] = layer_0[4351-:16] + bias_0[4351-:16];
                next_layer_0[4367-:16] = layer_0[4367-:16] + bias_0[4367-:16];
                next_layer_0[4383-:16] = layer_0[4383-:16] + bias_0[4383-:16];
                next_layer_0[4399-:16] = layer_0[4399-:16] + bias_0[4399-:16];
                next_layer_0[4415-:16] = layer_0[4415-:16] + bias_0[4415-:16];
                next_layer_0[4431-:16] = layer_0[4431-:16] + bias_0[4431-:16];
                next_layer_0[4447-:16] = layer_0[4447-:16] + bias_0[4447-:16];
                next_layer_0[4463-:16] = layer_0[4463-:16] + bias_0[4463-:16];
                next_layer_0[4479-:16] = layer_0[4479-:16] + bias_0[4479-:16];
                next_layer_0[4495-:16] = layer_0[4495-:16] + bias_0[4495-:16];
                next_layer_0[4511-:16] = layer_0[4511-:16] + bias_0[4511-:16];
                next_layer_0[4527-:16] = layer_0[4527-:16] + bias_0[4527-:16];
                next_layer_0[4543-:16] = layer_0[4543-:16] + bias_0[4543-:16];
                next_layer_0[4559-:16] = layer_0[4559-:16] + bias_0[4559-:16];
                next_layer_0[4575-:16] = layer_0[4575-:16] + bias_0[4575-:16];
                next_layer_0[4591-:16] = layer_0[4591-:16] + bias_0[4591-:16];
                next_layer_0[4607-:16] = layer_0[4607-:16] + bias_0[4607-:16];
                next_layer_0[4623-:16] = layer_0[4623-:16] + bias_0[4623-:16];
                next_layer_0[4639-:16] = layer_0[4639-:16] + bias_0[4639-:16];
                next_layer_0[4655-:16] = layer_0[4655-:16] + bias_0[4655-:16];
                next_layer_0[4671-:16] = layer_0[4671-:16] + bias_0[4671-:16];
                next_layer_0[4687-:16] = layer_0[4687-:16] + bias_0[4687-:16];
                next_layer_0[4703-:16] = layer_0[4703-:16] + bias_0[4703-:16];
                next_layer_0[4719-:16] = layer_0[4719-:16] + bias_0[4719-:16];
                next_layer_0[4735-:16] = layer_0[4735-:16] + bias_0[4735-:16];
                next_layer_0[4751-:16] = layer_0[4751-:16] + bias_0[4751-:16];
                next_layer_0[4767-:16] = layer_0[4767-:16] + bias_0[4767-:16];
                next_layer_0[4783-:16] = layer_0[4783-:16] + bias_0[4783-:16];
                next_layer_0[4799-:16] = layer_0[4799-:16] + bias_0[4799-:16];
                next_layer_0[4815-:16] = layer_0[4815-:16] + bias_0[4815-:16];
                next_layer_0[4831-:16] = layer_0[4831-:16] + bias_0[4831-:16];
                next_layer_0[4847-:16] = layer_0[4847-:16] + bias_0[4847-:16];
                next_layer_0[4863-:16] = layer_0[4863-:16] + bias_0[4863-:16];
                next_layer_0[4879-:16] = layer_0[4879-:16] + bias_0[4879-:16];
                next_layer_0[4895-:16] = layer_0[4895-:16] + bias_0[4895-:16];
                next_layer_0[4911-:16] = layer_0[4911-:16] + bias_0[4911-:16];
                next_layer_0[4927-:16] = layer_0[4927-:16] + bias_0[4927-:16];
                next_layer_0[4943-:16] = layer_0[4943-:16] + bias_0[4943-:16];
                next_layer_0[4959-:16] = layer_0[4959-:16] + bias_0[4959-:16];
                next_layer_0[4975-:16] = layer_0[4975-:16] + bias_0[4975-:16];
                next_layer_0[4991-:16] = layer_0[4991-:16] + bias_0[4991-:16];
                next_layer_0[5007-:16] = layer_0[5007-:16] + bias_0[5007-:16];
                next_layer_0[5023-:16] = layer_0[5023-:16] + bias_0[5023-:16];
                next_layer_0[5039-:16] = layer_0[5039-:16] + bias_0[5039-:16];
                next_layer_0[5055-:16] = layer_0[5055-:16] + bias_0[5055-:16];
                next_layer_0[5071-:16] = layer_0[5071-:16] + bias_0[5071-:16];
                next_layer_0[5087-:16] = layer_0[5087-:16] + bias_0[5087-:16];
                next_layer_0[5103-:16] = layer_0[5103-:16] + bias_0[5103-:16];
                next_layer_0[5119-:16] = layer_0[5119-:16] + bias_0[5119-:16];
                next_layer_0[5135-:16] = layer_0[5135-:16] + bias_0[5135-:16];
                next_layer_0[5151-:16] = layer_0[5151-:16] + bias_0[5151-:16];
                next_layer_0[5167-:16] = layer_0[5167-:16] + bias_0[5167-:16];
                next_layer_0[5183-:16] = layer_0[5183-:16] + bias_0[5183-:16];
                next_layer_0[5199-:16] = layer_0[5199-:16] + bias_0[5199-:16];
                next_layer_0[5215-:16] = layer_0[5215-:16] + bias_0[5215-:16];
                next_layer_0[5231-:16] = layer_0[5231-:16] + bias_0[5231-:16];
                next_layer_0[5247-:16] = layer_0[5247-:16] + bias_0[5247-:16];
                next_layer_0[5263-:16] = layer_0[5263-:16] + bias_0[5263-:16];
                next_layer_0[5279-:16] = layer_0[5279-:16] + bias_0[5279-:16];
                next_layer_0[5295-:16] = layer_0[5295-:16] + bias_0[5295-:16];
                next_layer_0[5311-:16] = layer_0[5311-:16] + bias_0[5311-:16];
                next_layer_0[5327-:16] = layer_0[5327-:16] + bias_0[5327-:16];
                next_layer_0[5343-:16] = layer_0[5343-:16] + bias_0[5343-:16];
                next_layer_0[5359-:16] = layer_0[5359-:16] + bias_0[5359-:16];
                next_layer_0[5375-:16] = layer_0[5375-:16] + bias_0[5375-:16];
                next_layer_0[5391-:16] = layer_0[5391-:16] + bias_0[5391-:16];
                next_layer_0[5407-:16] = layer_0[5407-:16] + bias_0[5407-:16];
                next_layer_0[5423-:16] = layer_0[5423-:16] + bias_0[5423-:16];
                next_layer_0[5439-:16] = layer_0[5439-:16] + bias_0[5439-:16];
                next_layer_0[5455-:16] = layer_0[5455-:16] + bias_0[5455-:16];
                next_layer_0[5471-:16] = layer_0[5471-:16] + bias_0[5471-:16];
                next_layer_0[5487-:16] = layer_0[5487-:16] + bias_0[5487-:16];
                next_layer_0[5503-:16] = layer_0[5503-:16] + bias_0[5503-:16];
                next_layer_0[5519-:16] = layer_0[5519-:16] + bias_0[5519-:16];
                next_layer_0[5535-:16] = layer_0[5535-:16] + bias_0[5535-:16];
                next_layer_0[5551-:16] = layer_0[5551-:16] + bias_0[5551-:16];
                next_layer_0[5567-:16] = layer_0[5567-:16] + bias_0[5567-:16];
                next_layer_0[5583-:16] = layer_0[5583-:16] + bias_0[5583-:16];
                next_layer_0[5599-:16] = layer_0[5599-:16] + bias_0[5599-:16];
                next_layer_0[5615-:16] = layer_0[5615-:16] + bias_0[5615-:16];
                next_layer_0[5631-:16] = layer_0[5631-:16] + bias_0[5631-:16];
                next_layer_0[5647-:16] = layer_0[5647-:16] + bias_0[5647-:16];
                next_layer_0[5663-:16] = layer_0[5663-:16] + bias_0[5663-:16];
                next_layer_0[5679-:16] = layer_0[5679-:16] + bias_0[5679-:16];
                next_layer_0[5695-:16] = layer_0[5695-:16] + bias_0[5695-:16];
                next_layer_0[5711-:16] = layer_0[5711-:16] + bias_0[5711-:16];
                next_layer_0[5727-:16] = layer_0[5727-:16] + bias_0[5727-:16];
                next_layer_0[5743-:16] = layer_0[5743-:16] + bias_0[5743-:16];
                next_layer_0[5759-:16] = layer_0[5759-:16] + bias_0[5759-:16];
                next_layer_0[5775-:16] = layer_0[5775-:16] + bias_0[5775-:16];
                next_layer_0[5791-:16] = layer_0[5791-:16] + bias_0[5791-:16];
                next_layer_0[5807-:16] = layer_0[5807-:16] + bias_0[5807-:16];
                next_layer_0[5823-:16] = layer_0[5823-:16] + bias_0[5823-:16];
                next_layer_0[5839-:16] = layer_0[5839-:16] + bias_0[5839-:16];
                next_layer_0[5855-:16] = layer_0[5855-:16] + bias_0[5855-:16];
                next_layer_0[5871-:16] = layer_0[5871-:16] + bias_0[5871-:16];
                next_layer_0[5887-:16] = layer_0[5887-:16] + bias_0[5887-:16];
                next_layer_0[5903-:16] = layer_0[5903-:16] + bias_0[5903-:16];
                next_layer_0[5919-:16] = layer_0[5919-:16] + bias_0[5919-:16];
                next_layer_0[5935-:16] = layer_0[5935-:16] + bias_0[5935-:16];
                next_layer_0[5951-:16] = layer_0[5951-:16] + bias_0[5951-:16];
                next_layer_0[5967-:16] = layer_0[5967-:16] + bias_0[5967-:16];
                next_layer_0[5983-:16] = layer_0[5983-:16] + bias_0[5983-:16];
                next_layer_0[5999-:16] = layer_0[5999-:16] + bias_0[5999-:16];
                next_layer_0[6015-:16] = layer_0[6015-:16] + bias_0[6015-:16];
                next_layer_0[6031-:16] = layer_0[6031-:16] + bias_0[6031-:16];
                next_layer_0[6047-:16] = layer_0[6047-:16] + bias_0[6047-:16];
                next_layer_0[6063-:16] = layer_0[6063-:16] + bias_0[6063-:16];
                next_layer_0[6079-:16] = layer_0[6079-:16] + bias_0[6079-:16];
                next_layer_0[6095-:16] = layer_0[6095-:16] + bias_0[6095-:16];
                next_layer_0[6111-:16] = layer_0[6111-:16] + bias_0[6111-:16];
                next_layer_0[6127-:16] = layer_0[6127-:16] + bias_0[6127-:16];
                next_layer_0[6143-:16] = layer_0[6143-:16] + bias_0[6143-:16];
                next_layer_0[6159-:16] = layer_0[6159-:16] + bias_0[6159-:16];
                next_layer_0[6175-:16] = layer_0[6175-:16] + bias_0[6175-:16];
                next_layer_0[6191-:16] = layer_0[6191-:16] + bias_0[6191-:16];
                next_layer_0[6207-:16] = layer_0[6207-:16] + bias_0[6207-:16];
                next_layer_0[6223-:16] = layer_0[6223-:16] + bias_0[6223-:16];
                next_layer_0[6239-:16] = layer_0[6239-:16] + bias_0[6239-:16];
                next_layer_0[6255-:16] = layer_0[6255-:16] + bias_0[6255-:16];
                next_layer_0[6271-:16] = layer_0[6271-:16] + bias_0[6271-:16];
                next_layer_0[6287-:16] = layer_0[6287-:16] + bias_0[6287-:16];
                next_layer_0[6303-:16] = layer_0[6303-:16] + bias_0[6303-:16];
                next_layer_0[6319-:16] = layer_0[6319-:16] + bias_0[6319-:16];
                next_layer_0[6335-:16] = layer_0[6335-:16] + bias_0[6335-:16];
                next_layer_0[6351-:16] = layer_0[6351-:16] + bias_0[6351-:16];
                next_layer_0[6367-:16] = layer_0[6367-:16] + bias_0[6367-:16];
                next_layer_0[6383-:16] = layer_0[6383-:16] + bias_0[6383-:16];
                next_layer_0[6399-:16] = layer_0[6399-:16] + bias_0[6399-:16];
                next_layer_0[6415-:16] = layer_0[6415-:16] + bias_0[6415-:16];
                next_layer_0[6431-:16] = layer_0[6431-:16] + bias_0[6431-:16];
                next_layer_0[6447-:16] = layer_0[6447-:16] + bias_0[6447-:16];
                next_layer_0[6463-:16] = layer_0[6463-:16] + bias_0[6463-:16];
                next_layer_0[6479-:16] = layer_0[6479-:16] + bias_0[6479-:16];
                next_layer_0[6495-:16] = layer_0[6495-:16] + bias_0[6495-:16];
                next_layer_0[6511-:16] = layer_0[6511-:16] + bias_0[6511-:16];
                next_layer_0[6527-:16] = layer_0[6527-:16] + bias_0[6527-:16];
                next_layer_0[6543-:16] = layer_0[6543-:16] + bias_0[6543-:16];
                next_layer_0[6559-:16] = layer_0[6559-:16] + bias_0[6559-:16];
                next_layer_0[6575-:16] = layer_0[6575-:16] + bias_0[6575-:16];
                next_layer_0[6591-:16] = layer_0[6591-:16] + bias_0[6591-:16];
                next_layer_0[6607-:16] = layer_0[6607-:16] + bias_0[6607-:16];
                next_layer_0[6623-:16] = layer_0[6623-:16] + bias_0[6623-:16];
                next_layer_0[6639-:16] = layer_0[6639-:16] + bias_0[6639-:16];
                next_layer_0[6655-:16] = layer_0[6655-:16] + bias_0[6655-:16];
                next_layer_0[6671-:16] = layer_0[6671-:16] + bias_0[6671-:16];
                next_layer_0[6687-:16] = layer_0[6687-:16] + bias_0[6687-:16];
                next_layer_0[6703-:16] = layer_0[6703-:16] + bias_0[6703-:16];
                next_layer_0[6719-:16] = layer_0[6719-:16] + bias_0[6719-:16];
                next_layer_0[6735-:16] = layer_0[6735-:16] + bias_0[6735-:16];
                next_layer_0[6751-:16] = layer_0[6751-:16] + bias_0[6751-:16];
                next_layer_0[6767-:16] = layer_0[6767-:16] + bias_0[6767-:16];
                next_layer_0[6783-:16] = layer_0[6783-:16] + bias_0[6783-:16];
                next_layer_0[6799-:16] = layer_0[6799-:16] + bias_0[6799-:16];
                next_layer_0[6815-:16] = layer_0[6815-:16] + bias_0[6815-:16];
                next_layer_0[6831-:16] = layer_0[6831-:16] + bias_0[6831-:16];
                next_layer_0[6847-:16] = layer_0[6847-:16] + bias_0[6847-:16];
                next_layer_0[6863-:16] = layer_0[6863-:16] + bias_0[6863-:16];
                next_layer_0[6879-:16] = layer_0[6879-:16] + bias_0[6879-:16];
                next_layer_0[6895-:16] = layer_0[6895-:16] + bias_0[6895-:16];
                next_layer_0[6911-:16] = layer_0[6911-:16] + bias_0[6911-:16];
                next_layer_0[6927-:16] = layer_0[6927-:16] + bias_0[6927-:16];
                next_layer_0[6943-:16] = layer_0[6943-:16] + bias_0[6943-:16];
                next_layer_0[6959-:16] = layer_0[6959-:16] + bias_0[6959-:16];
                next_layer_0[6975-:16] = layer_0[6975-:16] + bias_0[6975-:16];
                next_layer_0[6991-:16] = layer_0[6991-:16] + bias_0[6991-:16];
                next_layer_0[7007-:16] = layer_0[7007-:16] + bias_0[7007-:16];
                next_layer_0[7023-:16] = layer_0[7023-:16] + bias_0[7023-:16];
                next_layer_0[7039-:16] = layer_0[7039-:16] + bias_0[7039-:16];
                next_layer_0[7055-:16] = layer_0[7055-:16] + bias_0[7055-:16];
                next_layer_0[7071-:16] = layer_0[7071-:16] + bias_0[7071-:16];
                next_layer_0[7087-:16] = layer_0[7087-:16] + bias_0[7087-:16];
                next_layer_0[7103-:16] = layer_0[7103-:16] + bias_0[7103-:16];
                next_layer_0[7119-:16] = layer_0[7119-:16] + bias_0[7119-:16];
                next_layer_0[7135-:16] = layer_0[7135-:16] + bias_0[7135-:16];
                next_layer_0[7151-:16] = layer_0[7151-:16] + bias_0[7151-:16];
                next_layer_0[7167-:16] = layer_0[7167-:16] + bias_0[7167-:16];
                next_layer_0[7183-:16] = layer_0[7183-:16] + bias_0[7183-:16];
                next_layer_0[7199-:16] = layer_0[7199-:16] + bias_0[7199-:16];
                next_layer_0[7215-:16] = layer_0[7215-:16] + bias_0[7215-:16];
                next_layer_0[7231-:16] = layer_0[7231-:16] + bias_0[7231-:16];
                next_layer_0[7247-:16] = layer_0[7247-:16] + bias_0[7247-:16];
                next_layer_0[7263-:16] = layer_0[7263-:16] + bias_0[7263-:16];
                next_layer_0[7279-:16] = layer_0[7279-:16] + bias_0[7279-:16];
                next_layer_0[7295-:16] = layer_0[7295-:16] + bias_0[7295-:16];
                next_layer_0[7311-:16] = layer_0[7311-:16] + bias_0[7311-:16];
                next_layer_0[7327-:16] = layer_0[7327-:16] + bias_0[7327-:16];
                next_layer_0[7343-:16] = layer_0[7343-:16] + bias_0[7343-:16];
                next_layer_0[7359-:16] = layer_0[7359-:16] + bias_0[7359-:16];
                next_layer_0[7375-:16] = layer_0[7375-:16] + bias_0[7375-:16];
                next_layer_0[7391-:16] = layer_0[7391-:16] + bias_0[7391-:16];
                next_layer_0[7407-:16] = layer_0[7407-:16] + bias_0[7407-:16];
                next_layer_0[7423-:16] = layer_0[7423-:16] + bias_0[7423-:16];
                next_layer_0[7439-:16] = layer_0[7439-:16] + bias_0[7439-:16];
                next_layer_0[7455-:16] = layer_0[7455-:16] + bias_0[7455-:16];
                next_layer_0[7471-:16] = layer_0[7471-:16] + bias_0[7471-:16];
                next_layer_0[7487-:16] = layer_0[7487-:16] + bias_0[7487-:16];
                next_layer_0[7503-:16] = layer_0[7503-:16] + bias_0[7503-:16];
                next_layer_0[7519-:16] = layer_0[7519-:16] + bias_0[7519-:16];
                next_layer_0[7535-:16] = layer_0[7535-:16] + bias_0[7535-:16];
                next_layer_0[7551-:16] = layer_0[7551-:16] + bias_0[7551-:16];
                next_layer_0[7567-:16] = layer_0[7567-:16] + bias_0[7567-:16];
                next_layer_0[7583-:16] = layer_0[7583-:16] + bias_0[7583-:16];
                next_layer_0[7599-:16] = layer_0[7599-:16] + bias_0[7599-:16];
                next_layer_0[7615-:16] = layer_0[7615-:16] + bias_0[7615-:16];
                next_layer_0[7631-:16] = layer_0[7631-:16] + bias_0[7631-:16];
                next_layer_0[7647-:16] = layer_0[7647-:16] + bias_0[7647-:16];
                next_layer_0[7663-:16] = layer_0[7663-:16] + bias_0[7663-:16];
                next_layer_0[7679-:16] = layer_0[7679-:16] + bias_0[7679-:16];
                next_layer_0[7695-:16] = layer_0[7695-:16] + bias_0[7695-:16];
                next_layer_0[7711-:16] = layer_0[7711-:16] + bias_0[7711-:16];
                next_layer_0[7727-:16] = layer_0[7727-:16] + bias_0[7727-:16];
                next_layer_0[7743-:16] = layer_0[7743-:16] + bias_0[7743-:16];
                next_layer_0[7759-:16] = layer_0[7759-:16] + bias_0[7759-:16];
                next_layer_0[7775-:16] = layer_0[7775-:16] + bias_0[7775-:16];
                next_layer_0[7791-:16] = layer_0[7791-:16] + bias_0[7791-:16];
                next_layer_0[7807-:16] = layer_0[7807-:16] + bias_0[7807-:16];
                next_layer_0[7823-:16] = layer_0[7823-:16] + bias_0[7823-:16];
                next_layer_0[7839-:16] = layer_0[7839-:16] + bias_0[7839-:16];
                next_layer_0[7855-:16] = layer_0[7855-:16] + bias_0[7855-:16];
                next_layer_0[7871-:16] = layer_0[7871-:16] + bias_0[7871-:16];
                next_layer_0[7887-:16] = layer_0[7887-:16] + bias_0[7887-:16];
                next_layer_0[7903-:16] = layer_0[7903-:16] + bias_0[7903-:16];
                next_layer_0[7919-:16] = layer_0[7919-:16] + bias_0[7919-:16];
                next_layer_0[7935-:16] = layer_0[7935-:16] + bias_0[7935-:16];
                next_layer_0[7951-:16] = layer_0[7951-:16] + bias_0[7951-:16];
                next_layer_0[7967-:16] = layer_0[7967-:16] + bias_0[7967-:16];
                next_layer_0[7983-:16] = layer_0[7983-:16] + bias_0[7983-:16];
                next_layer_0[7999-:16] = layer_0[7999-:16] + bias_0[7999-:16];
                next_layer_0[8015-:16] = layer_0[8015-:16] + bias_0[8015-:16];
                next_layer_0[8031-:16] = layer_0[8031-:16] + bias_0[8031-:16];
                next_layer_0[8047-:16] = layer_0[8047-:16] + bias_0[8047-:16];
                next_layer_0[8063-:16] = layer_0[8063-:16] + bias_0[8063-:16];
                next_layer_0[8079-:16] = layer_0[8079-:16] + bias_0[8079-:16];
                next_layer_0[8095-:16] = layer_0[8095-:16] + bias_0[8095-:16];
                next_layer_0[8111-:16] = layer_0[8111-:16] + bias_0[8111-:16];
                next_layer_0[8127-:16] = layer_0[8127-:16] + bias_0[8127-:16];
                next_layer_0[8143-:16] = layer_0[8143-:16] + bias_0[8143-:16];
                next_layer_0[8159-:16] = layer_0[8159-:16] + bias_0[8159-:16];
                next_layer_0[8175-:16] = layer_0[8175-:16] + bias_0[8175-:16];
                next_layer_0[8191-:16] = layer_0[8191-:16] + bias_0[8191-:16];
                next_layer_0[8207-:16] = layer_0[8207-:16] + bias_0[8207-:16];
                next_layer_0[8223-:16] = layer_0[8223-:16] + bias_0[8223-:16];
                next_layer_0[8239-:16] = layer_0[8239-:16] + bias_0[8239-:16];
                next_layer_0[8255-:16] = layer_0[8255-:16] + bias_0[8255-:16];
                next_layer_0[8271-:16] = layer_0[8271-:16] + bias_0[8271-:16];
                next_layer_0[8287-:16] = layer_0[8287-:16] + bias_0[8287-:16];
                next_layer_0[8303-:16] = layer_0[8303-:16] + bias_0[8303-:16];
                next_layer_0[8319-:16] = layer_0[8319-:16] + bias_0[8319-:16];
                next_layer_0[8335-:16] = layer_0[8335-:16] + bias_0[8335-:16];
                next_layer_0[8351-:16] = layer_0[8351-:16] + bias_0[8351-:16];
                next_layer_0[8367-:16] = layer_0[8367-:16] + bias_0[8367-:16];
                next_layer_0[8383-:16] = layer_0[8383-:16] + bias_0[8383-:16];
                next_layer_0[8399-:16] = layer_0[8399-:16] + bias_0[8399-:16];
                next_layer_0[8415-:16] = layer_0[8415-:16] + bias_0[8415-:16];
                next_layer_0[8431-:16] = layer_0[8431-:16] + bias_0[8431-:16];
                next_layer_0[8447-:16] = layer_0[8447-:16] + bias_0[8447-:16];
                next_layer_0[8463-:16] = layer_0[8463-:16] + bias_0[8463-:16];
                next_layer_0[8479-:16] = layer_0[8479-:16] + bias_0[8479-:16];
                next_layer_0[8495-:16] = layer_0[8495-:16] + bias_0[8495-:16];
                next_layer_0[8511-:16] = layer_0[8511-:16] + bias_0[8511-:16];
                next_layer_0[8527-:16] = layer_0[8527-:16] + bias_0[8527-:16];
                next_layer_0[8543-:16] = layer_0[8543-:16] + bias_0[8543-:16];
                next_layer_0[8559-:16] = layer_0[8559-:16] + bias_0[8559-:16];
                next_layer_0[8575-:16] = layer_0[8575-:16] + bias_0[8575-:16];
                next_layer_0[8591-:16] = layer_0[8591-:16] + bias_0[8591-:16];
                next_layer_0[8607-:16] = layer_0[8607-:16] + bias_0[8607-:16];
                next_layer_0[8623-:16] = layer_0[8623-:16] + bias_0[8623-:16];
                next_layer_0[8639-:16] = layer_0[8639-:16] + bias_0[8639-:16];
                next_layer_0[8655-:16] = layer_0[8655-:16] + bias_0[8655-:16];
                next_layer_0[8671-:16] = layer_0[8671-:16] + bias_0[8671-:16];
                next_layer_0[8687-:16] = layer_0[8687-:16] + bias_0[8687-:16];
                next_layer_0[8703-:16] = layer_0[8703-:16] + bias_0[8703-:16];
                next_layer_0[8719-:16] = layer_0[8719-:16] + bias_0[8719-:16];
                next_layer_0[8735-:16] = layer_0[8735-:16] + bias_0[8735-:16];
                next_layer_0[8751-:16] = layer_0[8751-:16] + bias_0[8751-:16];
                next_layer_0[8767-:16] = layer_0[8767-:16] + bias_0[8767-:16];
                next_layer_0[8783-:16] = layer_0[8783-:16] + bias_0[8783-:16];
                next_layer_0[8799-:16] = layer_0[8799-:16] + bias_0[8799-:16];
                next_layer_0[8815-:16] = layer_0[8815-:16] + bias_0[8815-:16];
                next_layer_0[8831-:16] = layer_0[8831-:16] + bias_0[8831-:16];
                next_layer_0[8847-:16] = layer_0[8847-:16] + bias_0[8847-:16];
                next_layer_0[8863-:16] = layer_0[8863-:16] + bias_0[8863-:16];
                next_layer_0[8879-:16] = layer_0[8879-:16] + bias_0[8879-:16];
                next_layer_0[8895-:16] = layer_0[8895-:16] + bias_0[8895-:16];
                next_layer_0[8911-:16] = layer_0[8911-:16] + bias_0[8911-:16];
                next_layer_0[8927-:16] = layer_0[8927-:16] + bias_0[8927-:16];
                next_layer_0[8943-:16] = layer_0[8943-:16] + bias_0[8943-:16];
                next_layer_0[8959-:16] = layer_0[8959-:16] + bias_0[8959-:16];
                next_layer_0[8975-:16] = layer_0[8975-:16] + bias_0[8975-:16];
                next_layer_0[8991-:16] = layer_0[8991-:16] + bias_0[8991-:16];
                next_layer_0[9007-:16] = layer_0[9007-:16] + bias_0[9007-:16];
                next_layer_0[9023-:16] = layer_0[9023-:16] + bias_0[9023-:16];
                next_layer_0[9039-:16] = layer_0[9039-:16] + bias_0[9039-:16];
                next_layer_0[9055-:16] = layer_0[9055-:16] + bias_0[9055-:16];
                next_layer_0[9071-:16] = layer_0[9071-:16] + bias_0[9071-:16];
                next_layer_0[9087-:16] = layer_0[9087-:16] + bias_0[9087-:16];
                next_layer_0[9103-:16] = layer_0[9103-:16] + bias_0[9103-:16];
                next_layer_0[9119-:16] = layer_0[9119-:16] + bias_0[9119-:16];
                next_layer_0[9135-:16] = layer_0[9135-:16] + bias_0[9135-:16];
                next_layer_0[9151-:16] = layer_0[9151-:16] + bias_0[9151-:16];
                next_layer_0[9167-:16] = layer_0[9167-:16] + bias_0[9167-:16];
                next_layer_0[9183-:16] = layer_0[9183-:16] + bias_0[9183-:16];
                next_layer_0[9199-:16] = layer_0[9199-:16] + bias_0[9199-:16];
                next_layer_0[9215-:16] = layer_0[9215-:16] + bias_0[9215-:16];
                next_layer_0[9231-:16] = layer_0[9231-:16] + bias_0[9231-:16];
                next_layer_0[9247-:16] = layer_0[9247-:16] + bias_0[9247-:16];
                next_layer_0[9263-:16] = layer_0[9263-:16] + bias_0[9263-:16];
                next_layer_0[9279-:16] = layer_0[9279-:16] + bias_0[9279-:16];
                next_layer_0[9295-:16] = layer_0[9295-:16] + bias_0[9295-:16];
                next_layer_0[9311-:16] = layer_0[9311-:16] + bias_0[9311-:16];
                next_layer_0[9327-:16] = layer_0[9327-:16] + bias_0[9327-:16];
                next_layer_0[9343-:16] = layer_0[9343-:16] + bias_0[9343-:16];
                next_layer_0[9359-:16] = layer_0[9359-:16] + bias_0[9359-:16];
                next_layer_0[9375-:16] = layer_0[9375-:16] + bias_0[9375-:16];
                next_layer_0[9391-:16] = layer_0[9391-:16] + bias_0[9391-:16];
                next_layer_0[9407-:16] = layer_0[9407-:16] + bias_0[9407-:16];
                next_layer_0[9423-:16] = layer_0[9423-:16] + bias_0[9423-:16];
                next_layer_0[9439-:16] = layer_0[9439-:16] + bias_0[9439-:16];
                next_layer_0[9455-:16] = layer_0[9455-:16] + bias_0[9455-:16];
                next_layer_0[9471-:16] = layer_0[9471-:16] + bias_0[9471-:16];
                next_layer_0[9487-:16] = layer_0[9487-:16] + bias_0[9487-:16];
                next_layer_0[9503-:16] = layer_0[9503-:16] + bias_0[9503-:16];
                next_layer_0[9519-:16] = layer_0[9519-:16] + bias_0[9519-:16];
                next_layer_0[9535-:16] = layer_0[9535-:16] + bias_0[9535-:16];
                next_layer_0[9551-:16] = layer_0[9551-:16] + bias_0[9551-:16];
                next_layer_0[9567-:16] = layer_0[9567-:16] + bias_0[9567-:16];
                next_layer_0[9583-:16] = layer_0[9583-:16] + bias_0[9583-:16];
                next_layer_0[9599-:16] = layer_0[9599-:16] + bias_0[9599-:16];
                next_layer_0[9615-:16] = layer_0[9615-:16] + bias_0[9615-:16];
                next_layer_0[9631-:16] = layer_0[9631-:16] + bias_0[9631-:16];
                next_layer_0[9647-:16] = layer_0[9647-:16] + bias_0[9647-:16];
                next_layer_0[9663-:16] = layer_0[9663-:16] + bias_0[9663-:16];
                next_layer_0[9679-:16] = layer_0[9679-:16] + bias_0[9679-:16];
                next_layer_0[9695-:16] = layer_0[9695-:16] + bias_0[9695-:16];
                next_layer_0[9711-:16] = layer_0[9711-:16] + bias_0[9711-:16];
                next_layer_0[9727-:16] = layer_0[9727-:16] + bias_0[9727-:16];
                next_layer_0[9743-:16] = layer_0[9743-:16] + bias_0[9743-:16];
                next_layer_0[9759-:16] = layer_0[9759-:16] + bias_0[9759-:16];
                next_layer_0[9775-:16] = layer_0[9775-:16] + bias_0[9775-:16];
                next_layer_0[9791-:16] = layer_0[9791-:16] + bias_0[9791-:16];
                next_layer_0[9807-:16] = layer_0[9807-:16] + bias_0[9807-:16];
                next_layer_0[9823-:16] = layer_0[9823-:16] + bias_0[9823-:16];
                next_layer_0[9839-:16] = layer_0[9839-:16] + bias_0[9839-:16];
                next_layer_0[9855-:16] = layer_0[9855-:16] + bias_0[9855-:16];
                next_layer_0[9871-:16] = layer_0[9871-:16] + bias_0[9871-:16];
                next_layer_0[9887-:16] = layer_0[9887-:16] + bias_0[9887-:16];
                next_layer_0[9903-:16] = layer_0[9903-:16] + bias_0[9903-:16];
                next_layer_0[9919-:16] = layer_0[9919-:16] + bias_0[9919-:16];
                next_layer_0[9935-:16] = layer_0[9935-:16] + bias_0[9935-:16];
                next_layer_0[9951-:16] = layer_0[9951-:16] + bias_0[9951-:16];
                next_layer_0[9967-:16] = layer_0[9967-:16] + bias_0[9967-:16];
                next_layer_0[9983-:16] = layer_0[9983-:16] + bias_0[9983-:16];
                next_layer_0[9999-:16] = layer_0[9999-:16] + bias_0[9999-:16];
                next_layer_0[10015-:16] = layer_0[10015-:16] + bias_0[10015-:16];
                next_layer_0[10031-:16] = layer_0[10031-:16] + bias_0[10031-:16];
                next_layer_0[10047-:16] = layer_0[10047-:16] + bias_0[10047-:16];
                next_layer_0[10063-:16] = layer_0[10063-:16] + bias_0[10063-:16];
                next_layer_0[10079-:16] = layer_0[10079-:16] + bias_0[10079-:16];
                next_layer_0[10095-:16] = layer_0[10095-:16] + bias_0[10095-:16];
                next_layer_0[10111-:16] = layer_0[10111-:16] + bias_0[10111-:16];
                next_layer_0[10127-:16] = layer_0[10127-:16] + bias_0[10127-:16];
                next_layer_0[10143-:16] = layer_0[10143-:16] + bias_0[10143-:16];
                next_layer_0[10159-:16] = layer_0[10159-:16] + bias_0[10159-:16];
                next_layer_0[10175-:16] = layer_0[10175-:16] + bias_0[10175-:16];
                next_layer_0[10191-:16] = layer_0[10191-:16] + bias_0[10191-:16];
                next_layer_0[10207-:16] = layer_0[10207-:16] + bias_0[10207-:16];
                next_layer_0[10223-:16] = layer_0[10223-:16] + bias_0[10223-:16];
                next_layer_0[10239-:16] = layer_0[10239-:16] + bias_0[10239-:16];
                next_layer_0[10255-:16] = layer_0[10255-:16] + bias_0[10255-:16];
                next_layer_0[10271-:16] = layer_0[10271-:16] + bias_0[10271-:16];
                next_layer_0[10287-:16] = layer_0[10287-:16] + bias_0[10287-:16];
                next_layer_0[10303-:16] = layer_0[10303-:16] + bias_0[10303-:16];
                next_layer_0[10319-:16] = layer_0[10319-:16] + bias_0[10319-:16];
                next_layer_0[10335-:16] = layer_0[10335-:16] + bias_0[10335-:16];
                next_layer_0[10351-:16] = layer_0[10351-:16] + bias_0[10351-:16];
                next_layer_0[10367-:16] = layer_0[10367-:16] + bias_0[10367-:16];
                next_layer_0[10383-:16] = layer_0[10383-:16] + bias_0[10383-:16];
                next_layer_0[10399-:16] = layer_0[10399-:16] + bias_0[10399-:16];
                next_layer_0[10415-:16] = layer_0[10415-:16] + bias_0[10415-:16];
                next_layer_0[10431-:16] = layer_0[10431-:16] + bias_0[10431-:16];
                next_layer_0[10447-:16] = layer_0[10447-:16] + bias_0[10447-:16];
                next_layer_0[10463-:16] = layer_0[10463-:16] + bias_0[10463-:16];
                next_layer_0[10479-:16] = layer_0[10479-:16] + bias_0[10479-:16];
                next_layer_0[10495-:16] = layer_0[10495-:16] + bias_0[10495-:16];
                next_layer_0[10511-:16] = layer_0[10511-:16] + bias_0[10511-:16];
                next_layer_0[10527-:16] = layer_0[10527-:16] + bias_0[10527-:16];
                next_layer_0[10543-:16] = layer_0[10543-:16] + bias_0[10543-:16];
                next_layer_0[10559-:16] = layer_0[10559-:16] + bias_0[10559-:16];
                next_layer_0[10575-:16] = layer_0[10575-:16] + bias_0[10575-:16];
                next_layer_0[10591-:16] = layer_0[10591-:16] + bias_0[10591-:16];
                next_layer_0[10607-:16] = layer_0[10607-:16] + bias_0[10607-:16];
                next_layer_0[10623-:16] = layer_0[10623-:16] + bias_0[10623-:16];
                next_layer_0[10639-:16] = layer_0[10639-:16] + bias_0[10639-:16];
                next_layer_0[10655-:16] = layer_0[10655-:16] + bias_0[10655-:16];
                next_layer_0[10671-:16] = layer_0[10671-:16] + bias_0[10671-:16];
                next_layer_0[10687-:16] = layer_0[10687-:16] + bias_0[10687-:16];
                next_layer_0[10703-:16] = layer_0[10703-:16] + bias_0[10703-:16];
                next_layer_0[10719-:16] = layer_0[10719-:16] + bias_0[10719-:16];
                next_layer_0[10735-:16] = layer_0[10735-:16] + bias_0[10735-:16];
                next_layer_0[10751-:16] = layer_0[10751-:16] + bias_0[10751-:16];
                next_layer_0[10767-:16] = layer_0[10767-:16] + bias_0[10767-:16];
                next_layer_0[10783-:16] = layer_0[10783-:16] + bias_0[10783-:16];
                next_layer_0[10799-:16] = layer_0[10799-:16] + bias_0[10799-:16];
                next_layer_0[10815-:16] = layer_0[10815-:16] + bias_0[10815-:16];
                next_layer_0[10831-:16] = layer_0[10831-:16] + bias_0[10831-:16];
                next_layer_0[10847-:16] = layer_0[10847-:16] + bias_0[10847-:16];
                next_layer_0[10863-:16] = layer_0[10863-:16] + bias_0[10863-:16];
                next_layer_0[10879-:16] = layer_0[10879-:16] + bias_0[10879-:16];
                next_layer_0[10895-:16] = layer_0[10895-:16] + bias_0[10895-:16];
                next_layer_0[10911-:16] = layer_0[10911-:16] + bias_0[10911-:16];
                next_layer_0[10927-:16] = layer_0[10927-:16] + bias_0[10927-:16];
                next_layer_0[10943-:16] = layer_0[10943-:16] + bias_0[10943-:16];
                next_layer_0[10959-:16] = layer_0[10959-:16] + bias_0[10959-:16];
                next_layer_0[10975-:16] = layer_0[10975-:16] + bias_0[10975-:16];
                next_layer_0[10991-:16] = layer_0[10991-:16] + bias_0[10991-:16];
                next_layer_0[11007-:16] = layer_0[11007-:16] + bias_0[11007-:16];
                next_layer_0[11023-:16] = layer_0[11023-:16] + bias_0[11023-:16];
                next_layer_0[11039-:16] = layer_0[11039-:16] + bias_0[11039-:16];
                next_layer_0[11055-:16] = layer_0[11055-:16] + bias_0[11055-:16];
                next_layer_0[11071-:16] = layer_0[11071-:16] + bias_0[11071-:16];
                next_layer_0[11087-:16] = layer_0[11087-:16] + bias_0[11087-:16];
                next_layer_0[11103-:16] = layer_0[11103-:16] + bias_0[11103-:16];
                next_layer_0[11119-:16] = layer_0[11119-:16] + bias_0[11119-:16];
                next_layer_0[11135-:16] = layer_0[11135-:16] + bias_0[11135-:16];
                next_layer_0[11151-:16] = layer_0[11151-:16] + bias_0[11151-:16];
                next_layer_0[11167-:16] = layer_0[11167-:16] + bias_0[11167-:16];
                next_layer_0[11183-:16] = layer_0[11183-:16] + bias_0[11183-:16];
                next_layer_0[11199-:16] = layer_0[11199-:16] + bias_0[11199-:16];
                next_layer_0[11215-:16] = layer_0[11215-:16] + bias_0[11215-:16];
                next_layer_0[11231-:16] = layer_0[11231-:16] + bias_0[11231-:16];
                next_layer_0[11247-:16] = layer_0[11247-:16] + bias_0[11247-:16];
                next_layer_0[11263-:16] = layer_0[11263-:16] + bias_0[11263-:16];
                next_layer_0[11279-:16] = layer_0[11279-:16] + bias_0[11279-:16];
                next_layer_0[11295-:16] = layer_0[11295-:16] + bias_0[11295-:16];
                next_layer_0[11311-:16] = layer_0[11311-:16] + bias_0[11311-:16];
                next_layer_0[11327-:16] = layer_0[11327-:16] + bias_0[11327-:16];
                next_layer_0[11343-:16] = layer_0[11343-:16] + bias_0[11343-:16];
                next_layer_0[11359-:16] = layer_0[11359-:16] + bias_0[11359-:16];
                next_layer_0[11375-:16] = layer_0[11375-:16] + bias_0[11375-:16];
                next_layer_0[11391-:16] = layer_0[11391-:16] + bias_0[11391-:16];
                next_layer_0[11407-:16] = layer_0[11407-:16] + bias_0[11407-:16];
                next_layer_0[11423-:16] = layer_0[11423-:16] + bias_0[11423-:16];
                next_layer_0[11439-:16] = layer_0[11439-:16] + bias_0[11439-:16];
                next_layer_0[11455-:16] = layer_0[11455-:16] + bias_0[11455-:16];
                next_layer_0[11471-:16] = layer_0[11471-:16] + bias_0[11471-:16];
                next_layer_0[11487-:16] = layer_0[11487-:16] + bias_0[11487-:16];
                next_layer_0[11503-:16] = layer_0[11503-:16] + bias_0[11503-:16];
                next_layer_0[11519-:16] = layer_0[11519-:16] + bias_0[11519-:16];
                next_layer_0[11535-:16] = layer_0[11535-:16] + bias_0[11535-:16];
                next_layer_0[11551-:16] = layer_0[11551-:16] + bias_0[11551-:16];
                next_layer_0[11567-:16] = layer_0[11567-:16] + bias_0[11567-:16];
                next_layer_0[11583-:16] = layer_0[11583-:16] + bias_0[11583-:16];
                next_layer_0[11599-:16] = layer_0[11599-:16] + bias_0[11599-:16];
                next_layer_0[11615-:16] = layer_0[11615-:16] + bias_0[11615-:16];
                next_layer_0[11631-:16] = layer_0[11631-:16] + bias_0[11631-:16];
                next_layer_0[11647-:16] = layer_0[11647-:16] + bias_0[11647-:16];
                next_layer_0[11663-:16] = layer_0[11663-:16] + bias_0[11663-:16];
                next_layer_0[11679-:16] = layer_0[11679-:16] + bias_0[11679-:16];
                next_layer_0[11695-:16] = layer_0[11695-:16] + bias_0[11695-:16];
                next_layer_0[11711-:16] = layer_0[11711-:16] + bias_0[11711-:16];
                next_layer_0[11727-:16] = layer_0[11727-:16] + bias_0[11727-:16];
                next_layer_0[11743-:16] = layer_0[11743-:16] + bias_0[11743-:16];
                next_layer_0[11759-:16] = layer_0[11759-:16] + bias_0[11759-:16];
                next_layer_0[11775-:16] = layer_0[11775-:16] + bias_0[11775-:16];
                next_layer_0[11791-:16] = layer_0[11791-:16] + bias_0[11791-:16];
                next_layer_0[11807-:16] = layer_0[11807-:16] + bias_0[11807-:16];
                next_layer_0[11823-:16] = layer_0[11823-:16] + bias_0[11823-:16];
                next_layer_0[11839-:16] = layer_0[11839-:16] + bias_0[11839-:16];
                next_layer_0[11855-:16] = layer_0[11855-:16] + bias_0[11855-:16];
                next_layer_0[11871-:16] = layer_0[11871-:16] + bias_0[11871-:16];
                next_layer_0[11887-:16] = layer_0[11887-:16] + bias_0[11887-:16];
                next_layer_0[11903-:16] = layer_0[11903-:16] + bias_0[11903-:16];
                next_layer_0[11919-:16] = layer_0[11919-:16] + bias_0[11919-:16];
                next_layer_0[11935-:16] = layer_0[11935-:16] + bias_0[11935-:16];
                next_layer_0[11951-:16] = layer_0[11951-:16] + bias_0[11951-:16];
                next_layer_0[11967-:16] = layer_0[11967-:16] + bias_0[11967-:16];
                next_layer_0[11983-:16] = layer_0[11983-:16] + bias_0[11983-:16];
                next_layer_0[11999-:16] = layer_0[11999-:16] + bias_0[11999-:16];
                next_layer_0[12015-:16] = layer_0[12015-:16] + bias_0[12015-:16];
                next_layer_0[12031-:16] = layer_0[12031-:16] + bias_0[12031-:16];
                next_layer_0[12047-:16] = layer_0[12047-:16] + bias_0[12047-:16];
                next_layer_0[12063-:16] = layer_0[12063-:16] + bias_0[12063-:16];
                next_layer_0[12079-:16] = layer_0[12079-:16] + bias_0[12079-:16];
                next_layer_0[12095-:16] = layer_0[12095-:16] + bias_0[12095-:16];
                next_layer_0[12111-:16] = layer_0[12111-:16] + bias_0[12111-:16];
                next_layer_0[12127-:16] = layer_0[12127-:16] + bias_0[12127-:16];
                next_layer_0[12143-:16] = layer_0[12143-:16] + bias_0[12143-:16];
                next_layer_0[12159-:16] = layer_0[12159-:16] + bias_0[12159-:16];
                next_layer_0[12175-:16] = layer_0[12175-:16] + bias_0[12175-:16];
                next_layer_0[12191-:16] = layer_0[12191-:16] + bias_0[12191-:16];
                next_layer_0[12207-:16] = layer_0[12207-:16] + bias_0[12207-:16];
                next_layer_0[12223-:16] = layer_0[12223-:16] + bias_0[12223-:16];
                next_layer_0[12239-:16] = layer_0[12239-:16] + bias_0[12239-:16];
                next_layer_0[12255-:16] = layer_0[12255-:16] + bias_0[12255-:16];
                next_layer_0[12271-:16] = layer_0[12271-:16] + bias_0[12271-:16];
                next_layer_0[12287-:16] = layer_0[12287-:16] + bias_0[12287-:16];
                next_layer_0[12303-:16] = layer_0[12303-:16] + bias_0[12303-:16];
                next_layer_0[12319-:16] = layer_0[12319-:16] + bias_0[12319-:16];
                next_layer_0[12335-:16] = layer_0[12335-:16] + bias_0[12335-:16];
                next_layer_0[12351-:16] = layer_0[12351-:16] + bias_0[12351-:16];
                next_layer_0[12367-:16] = layer_0[12367-:16] + bias_0[12367-:16];
                next_layer_0[12383-:16] = layer_0[12383-:16] + bias_0[12383-:16];
                next_layer_0[12399-:16] = layer_0[12399-:16] + bias_0[12399-:16];
                next_layer_0[12415-:16] = layer_0[12415-:16] + bias_0[12415-:16];
                next_layer_0[12431-:16] = layer_0[12431-:16] + bias_0[12431-:16];
                next_layer_0[12447-:16] = layer_0[12447-:16] + bias_0[12447-:16];
                next_layer_0[12463-:16] = layer_0[12463-:16] + bias_0[12463-:16];
                next_layer_0[12479-:16] = layer_0[12479-:16] + bias_0[12479-:16];
                next_layer_0[12495-:16] = layer_0[12495-:16] + bias_0[12495-:16];
                next_layer_0[12511-:16] = layer_0[12511-:16] + bias_0[12511-:16];
                next_layer_0[12527-:16] = layer_0[12527-:16] + bias_0[12527-:16];
                next_layer_0[12543-:16] = layer_0[12543-:16] + bias_0[12543-:16];

            end
            SFIN: begin
                next_layer_0 = layer_0;
            end
            default: begin
                next_layer_0 = layer_0;
            end
        endcase
    end
endmodule